`timescale 1ns / 1ps
`include "../../sources_1/new/defines.v"
module lw_hmac_tb;
/*
  key_s32: 09a09c09c989a09023b432e28000323f87c79a9008f0ff323225656e3326234fca889df080bc09a3bc54d2af4b23c26e32bb2af423e2a24c4f5233c599c7689e
  key_s64: 07f089fd09a09c09890b9089c989a0904542345f23b432e2a98b09c98000323f089b977987c79a90b4c6ba9908f0ff32665253463225656e62546a453326234f9809b908ca889df06877a9d980bc09a343525245bc54d2af6c2345d34b23c26e624352e332bb2af44525232f23e2a24c253456324f5233c5a9877b9899c7689e
  simple_key_s32: 0000000c0000000d0000000a0000000b00000008000000090000009000000080000000f0000000e0000000d0000000c000000c0000000d0000000a0000000b0f
  simple_key_s64: 000000000000000c000000000000000d000000000000000a000000000000000b000000000000000800000000000000090000000000000090000000000000008000000000000000f000000000000000e000000000000000d000000000000000c00000000000000c000000000000000d000000000000000a000000000000000b0f

  test cases S32:
  test 1 - NULL
  test 2 - abc
  test 3 - abcdbcdecdefdefgefghfghighijhijkijkljklmklmnlmnomnopnopq
  test 4 - rewqiuytsapohgfd;lkjcxz'mbnvf/.,nbedxvium,aw5duinuerfxsbvbastyxmoiuytrewgfdslkjh,mnbvcxzxzaqwsxcedcvrfvbtgbnyhnmujm,rewqiuytsapohgfd;lkjcxz'mbnvf/.,
  test 5 - 88866d5a04c2b81f579962b7293928a6a2458381ef4f022fc2ec7a72422b275e0f5588e36c63f371a4ddd72d89308a6d1a41e5edced3f805720ecea64f09d21b1059ff90b5b1f5e9ff7f3374da3ded1d47eb9f6562d0bff48974c0234e5be5fa1f571c984c5d4dc8edbd13d4fffc20b5009578b782b7f6b029d1b1b4c7726ef8870d1b9130d967e6b170352e3c1d04579ad3f1207efca01c6d0d4416329e118a66fb0974bac9a026e5511650a4a2a1c10264cf24c38d0c66f3cf3102e2c5be3e69ffd24fcf964f94dcc329543f8be0b67d3ec91547a61ce928ff1e2d1072c1ab9b499dda9a37847747d0011f6457f03dafdce9e23ea6bbbf4371eae2b4278f914ac099c428bdac62d9e0e28a8c97dfd9942a26bb9323b199787ec001a4fc7d8cda3db0928947ddaa9c73dd1a5a496d6e86adaca8ef5b071bda3269f9a31629d8
  test 6 - d364e8f1545ce324431f92858db5d670dbb90c597149fd94402fbef07d04a3f76e5604c98102eec5adb391582c6758b85ddd03f53b1696b125c71235cf692dd45f260dd4fe1e19759544655511310ce88581166caa512601073ddceaa9a0d3608952ecd51bf2a12ed18ad3d8a246c2098d97d8dc762483c49ce8e1ccb4c7ff8721b765046af02a3b44fa8a4ffb474e3c8dfc121c7a4fcf5cf597b269b8465ed838be2884645a504f251846bd82e8ccdcc7f4296b6995d44fd2b3634322c119a11abdcff594756536f1d217d65dfcc6e48dfe4976865425f17f95f9b420368ea99df22598c33f49b0a9f669485e5661682d698fc973c0e1b4627d53fe417e82be13243d29ef5c950f56cb298cedbffac5899ca76c4e785cf683468eb897aca16e0438df074093b0e177e94d707ebece79fe133407a7f48756c5d112f3de2ff50e
  test 7 - 010010000111000001011110100110010100010011011010010001001011010011001000000100111000111100110000100000011010000000000001110100101111001010001010110011000001011001110100010101101011001011000111011110110011011001101011110011000001110010000001010001110100010111001100011000010001010011010111011010111100110001000010010000111000000110110101010001010011111011000111100000110011101101111101111010011100001011001111000011111000101000011000010111011110111110001000011110110101011111011010100000101010001011100111010111101001100010111001110101010011010001110010010110011010110011001111100001001011011100011000001101011001000000011100100100110000111001101100100101010100000011111010000001011110101100010111001010001010010011010101010000110010010101110000011011011100100011110001001101011110000101101001010110000110001101101011110010010111111101011010100000111101000010111110111001000101001101010000101011010000001101101011111010011000001011101110101101100010101010011010010101101010110011111000010101011110110111001010001101000010011100101001001111111001100011101100010001011110100111100010011111001000101001111111001101011000000011001100000100001011110010000100001101111010110010010000010011010100110001100001110111000110110000100110011010010011111100010011000000101010000101110001001010001111111000111101001010101001100000100001101110100011111111101110100111000001010100001110001001001111001110110001110110111000100011111100000011111110000000110010011111010011011101101100011110011100011100101101111000000111101101101101101011001000000110110011101101000010111001100000001111111110110010000010100011111100000110001010110000100101010100010111011010111100101111000111010010010100000011111111101101001101100001111111011000111111110100100100000100110000100111011101100000010001010111011000000100101000011010011011010110010101110101101110010011111010111001011100111010000111101010110100000010110000010010000111101111100001110111101100110000000010010011111101001101111011000110000001101101101001110010110100011000101110000110110001001011100100011110010000111100000000111111111011100011011100001110001011110110001101011100010111110000101000111010001100110101100000110101000001111011000001111111111100000100111100111110001110110010000010100110100011011001101100100111111011001111011101111000100011100100110011101101011000101011101100010100101110110001101010111110100110000101011100100001101010010110100010000011010101010011011100010111011111101101101111000110100011000000011001100011111000110010100111100101011011100101110010000011010101111010110011110001111000000111100100101110110010010001001100000111110111100011100010011100011101001000110001011111111000011000010001001111010100001011000011000000011011101100100010010110011101111110000011111001010000010001000011010111001000010111100100101001100110111111010111100010010010001011111011011011100100110101111010010010111011111011100110010110101110010101111101001110111110000000000101010011110111011101011010010010011010000101011100010100101010111011010101110110111100100010111011101000001110000110111110111111001011000101110011111110101011001010010100111111010000011111001001110101011110011101111101000010100110100001101010100000101001001001001000101000101001000110000011010111111110010001111010111110011010011001010001101010100100000010001101101010111010110101000100100111010110100011110001010010000101110000000101110011011101101110110111000110011101110000010000100000001000101110100000000011001110011110000110101100101011110100000010001110010111011000000100110010011110100100000111001101010001000100111110101101111011001011011110001110010000100100010010010110001111000011011101010001101010110110000011000010110001010010000010010111010100011000011001111100100110111110111011001010010111101101110001110100001011100100000000011111000000101010100101100011111001010010010011000110100001110010100001001001100001101100101111010110111100001001010101110001010011110001111101001000110000100001110101111110101101111011111001100101111001101011100
  
  test cases S64:
  test 1 - NULL
  test 2 - abc
  test 3 - abcdefghbcdefghicdefghijdefghijkefghijklfghijklmghijklmnhijklmnoijklmnopjklmnopqklmnopqrlmnopqrsmnopqrstnopqrstu
  test 4 - aaaarewqaaaaiuytaaaasapoaaaahgfdaaaa;lkjaaaacxz'aaaambnvaaaaf/.,aaaanbedaaaaxviuaaaam,awaaaa5duiaaaanueraaaafxsbaaaavbasaaaatyxmaaaaoiuyaaaatrewaaaagfdsaaaalkjhaaaa,mnbaaaavcxzaaaaxzaqaaaawsxcaaaaedcvaaaarfvbaaaatgbnaaaayhnmaaaaujm,aaaarewqaaaaiuytaaaasapoaaaahgfdaaaa;lkjaaaacxz'aaaambnvaaaaf/.,
  test 5 - e6e3f8e688866d5aace56b5104c2b81f2018c313579962b7c6354eca293928a653c3ce94a24583810a4d1749ef4f022fb650afa7c2ec7a727f45199c422b275e0c6676b60f5588e307bd2fe86c63f3712f161f70a4ddd72df9373e2d89308a6df583789d1a41e5edca6ad14eced3f8054d0644ba720ecea679fc057f4f09d21b49e657721059ff90c877faf0b5b1f5e9e0f4e816ff7f3374e41907aada3ded1da34aa42947eb9f651ad3757262d0bff41fca46548974c023a6b97ea34e5be5fa3123ee961f571c98c2163b7f4c5d4dc896c0163dedbd13d403feb51cfffc20b5924ff032009578b71094c54782b7f6b007f9687229d1b1b46fecd110c7726ef8deafb5db870d1b91a3dfecba30d967e624b722a3b170352ea50cb10d3c1d0457ebfc6f9a9ad3f1205daf2cbc7efca01c178bbd696d0d44163e214615329e118ac4f8f82d66fb0974255ec7a0bac9a026bfff2feee5511650aac079fba4a2a1c17c3dafdd0264cf241242500dc38d0c663e56ebc4f3cf31020fdce116e2c5be3ed9d590cb69ffd24f036cb56fcf964f94d4f5c702dcc32954f0dab7533f8be0b6eaae6e6e7d3ec915ec7f4a1347a61ce9af868f7528ff1e2d528add981072c1ab107a9c2f9b499dda34e11d2a9a37847780a2b49647d0011f63e7fd806457f03d5c33fa38afdce9e2fe6f618c3ea6bbbf4e54d9e04371eae2764c1ef7b4278f911027361f4ac099c4fa9d1e0028bdac622b669e27d9e0e28a3d93e0598c97dfd95fa61c62942a26bb2abf21e19323b19923442d99787ec0013f694bf9a4fc7d8cdcdd6339da3db0929af7b8e58947ddaac137331f9c73dd1aa9c62a685a496d6e9991e65286adaca8e9b8263eef5b071bcdaa1882da3269f90cebdb81a31629d8
  tset 6 - 7794cc3dd364e8f1e09d1a01545ce3245507945b431f92855bfc5e6c8db5d6703a70f2a4dbb90c59277e4d9b7149fd943e1f2098402fbef06e91e2bf7d04a3f7d52c59156e5604c9a00c386b8102eec58b4d7516adb391582a2631ae2c6758b8fa14ee1c5ddd03f500deb1fe3b1696b19bdc06a725c71235c19bf174cf692dd4873228985f260dd4df2a943afe1e1975a0376d409544655565e5752911310ce8bbaf26338581166c1ae70046aa512601f6f5cfc0073ddcea1e98d569a9a0d360f1852d1c8952ecd596e6bca81bf2a12e61e26ba9d18ad3d8a25aa131a246c209da976c748d97d8dcddce6ad5762483c463404bdf9ce8e1cc3aa29fe6b4c7ff87e6bf8a6821b76504ba61dea66af02a3b3ff028c444fa8a4f256333e6fb474e3c707b78758dfc121c9f38ecc97a4fcf5c8a0a9995f597b26944a54e5fb8465ed8f327255438be2884e0334b97645a504f42d7fd66251846bd8dfc70da82e8ccdc1ca860d2c7f4296b91353bae6995d44f4a7b69dad2b36343b0fca6e922c119a1ddd0f86d1abdcff5f47084e4947565361394f23af1d217d65342c6285dfcc6e4a39cc4928dfe4976b07d6156865425f1129438387f95f9b44718e6f720368ea9e51cb8289df2259899bb3a2cc33f49b0bde2c64ea9f66948bf9043885e566168a087ce262d698fc99b1eed3273c0e1b4dd477829627d53fe17c16b85417e82bee21ac93e13243d29b9b5cb46ef5c950f420d2c9656cb298c03913407edbffac57db4cbcd899ca76c7b8582b54e785cf692ab7be983468eb82784bbb497aca16e7bfd75590438df07e1c0e7874093b0e1fd73f25d77e94d70f823391d7ebece79f3a929cefe133407aa9cf54fa7f48756712c2ec4c5d112f380077bc3de2ff50e
  test 7 - 000010101011100001101111111101000100100001110000010111101001100110010100100101011001111101001101010001001101101001000100101101000001001111000000011011000011111011001000000100111000111100110000011101110011010101110000010011011000000110100000000000011101001000111100010011000011000100110101111100101000101011001100000101100100000100111110100101111000110101110100010101101011001011000111110110001110010110100100101001010111101100110110011010111100110000011001110000110101111110110001000111001000000101000111010001010111110101000110000100010010100111001100011000010001010011010111101010000100101010110100011011110110101111001100010000100100001110000101111000001010100110110011100000011011010101000101001111101001100001001110101010010001010011000111100000110011101101111101100100000101011111111110000001111110100111000010110011110000111100011100101111001111001111111101100010100001100001011101111011110000000000000010100010010100000010001000011110110101011111011010011010000111011001101011000111101000001010100010111001110101111001111100011011110010010001001010100110001011100111010101001101001010001101001101001110010000011101110010010110011010110011001111111101101110110111001001000001101000010010110111000110000011010101100011111000011100000000101011100100000001110010010011000011100010101110101000010110111111111101101100100101010100000011111010000110101010110001010001000100000000010111101011000101110010100010000111111100110011010000000100101001001101010101000011001001011101011111100000111001100010000001110000011011011100100011110001110000010000001100001011100100010011010111100001011010010101100000000010000011100011001101100001011000110110101111001001011111111001110001011111010100111101100001011010100000111101000010111110101100100001000011111010100001101110010001010011010100001010110101001000100101000010000011100111000000110110101111101001100000101110010111100011010001011100000011101110101101100010101010011010010110101001100100100101010110000101011010101100111110000101010100100111101101001000111100101000111011011100101000110100001001111100110111000000101011100011111000101001001111111001100011101100111001110011010110100111110100110100010111101001111000100111110010011000100001000011100010100000100010100111111100110101100000001010000000011010101010110011111111001100000100001011110010000100100110110101110001111111000011000011011110101100100100000100110110111110010110000010000111100110010011000110000111011100011011000001000000101101100001011001001100100110011010010011111100010011101100010010000000110000000100000000001010100001011100010010100001101010100010011110010101011101111111100011110100101010100110000110000101000000101101000100101100100001101110100011111111101110000011010111000100100111111101001001110000010101000011100010010010110101101011001010110100110001010011110011101100011101101110000111110111111011110110110110011110001111110000001111111000000011111110110111010001110010000001100010011111010011011101101100011110111011010100111111100111000000100111000111001011011110000001111010111001001101100110011110110010110110110110101100100000011011111001110101110010110001011110110011101101000010111001100000001110001111101110101111010001111101111111101100100000101000111111001101010111011011101010011101001000011000101011000010010101010001000010011111110101001001000101110111011010111100101111000111010000001011110010001011001110111101100101000000111111111011010011011011000101001110111111011000111010000111111101100011111111010010111001101110110000111101100010000100000100110000100111011101100010010001100100110100011100110011000100010101110110000001001010000010111011110111010110011100001001101001101101011001010111010110110111011100010111000010100100001110010011111010111001011100111010111111011000101100100101100110100001111010101101000000101100000100010010100101010011101111001001001000011110111110000111011110011011011100010110101111000000101100110000000010010011111101001111001110100100010010011011000001011101011011000110000001101101100011011011110001001111101011010010011100000010110100011000101110111100000110101110010111011001100001101100010010111001000111100101110010100100100101100111000000000011110000000011111111101110001100101010011101001111110011100111011100001110001011110110001101000110101011010000100001010111000111000101111100001010001110100010011001110001101000010010101001110011010110000011010100000111101001001001111011101111100010110011000001111111111100000100111100101100000110101101011011010101011111100011101100100000101001101001111000100011011100000000000011001101100110110010011111101100110001011111110010000011101110001011011101111000100011100100110011010111101011001101001001111101111011010110001010111011000101001010110010100010111010011110010100111011000110101011111010011000011010010110101001000111100011011101011100100001101010010110100010101110111011110011110100011100110000110101010100110111000101110101100001010101100011111001011000111110110110111100011010001100001100110000011001001111111100100100011001100011111000110010100111000000011001100111101110000000011001010110111001011100100000110101110010111110100000010011011011010111101011001111000111100000011011110000001011010111111011001011100100101110110010010001001100011001100011011000010111001010000001111101111000111000100111000111010000011000110000001000000111110100100011000101111111100001101010100110111001100110101001110000010001001111010100001011000011111100001111001010000111111000000000000110111011001000100101100110000111110011011101101100011100110111111000001111100101000001000000100111111100111100001000011101000011010111001000010111100100011010001100000101000101000010011010011001101111110101111000100110100000111001011111001110100011001000101111101101101110010011011011100011111110110011011110101101111010010010111011111011100110101000000100010000111100000111010101101011100101011111010011101111000001110111001111101010100111111000000000010101001111011101110110011001010101000101010101001001011010010010011010000101011100000010101001000001001111111100010101001010101110110101011101101111000000111100000111100110011010110010001011101110100000111000010010101111110111000000110100100110111110111111001011000101110011001011101010001111010010000100001111101010110010100101001111110110000000101110001110010101110011000001111100100111010101111001110001011011000001000100010110010101111101000010100110100001101010111011101100101111011100101001011000001010010010010010001010001001110000000111000011001100101111100100011000001101011111111001001111001011111001110000011100000101111010111110011010011001010001111001001000010100111001010001011010101001000000100011011010101111010110011101110100001111000110101011010100010010011101011010001011110011001011011111101011000111110001010010000101110000000101011000101110010001001100001101101100110111011011011100011001110101000111000110010011111111101110110000010000100000001000101110101010011100001100111011000001111100000000110011100111100001101011010010101001010011010000011100010010101111010000001000111001011111010111111100011100111011011011011000000100110010011110100100001011000100101010000111100001101001110011010100010001001111101011110011100010100001101100100100110111101100101101111000111001000001110101001111010100101111011100100100010010010110001111000011011100001010001011100101011100011011010100011010101101100000110000000110110111111110010001001100011011000101001000001001011101010001000101011100110000011010100101011000011001111100100110111110110110111101000110100011010111000110110010100101111011011100011101101111001000110000110111101101000000101110010000000001111100000010110100100100101101000001111001101010100101100011111001010010011001110001100010101011110101100100110001101000011100101000010010010101010110001101100110010010010110000110110010111101011011110010001100111011001000001100001111001001010101110001010011110001110010010110100000001010000001010011010010001100001000011101011111011101011100111101111101101101011010110111101111100110010111100111111010010100110000000001000011101011100
*/
  logic clk_i;
  logic aresetn_i;
  logic start_i;
  logic abort_i = 1'b0;
  logic last_i;
  logic data_valid_i;
  logic [`WORD_SIZE-1:0] data_i;
  logic [1:0] random_i;
  logic [3:0] opcode_i;
  logic [`WORD_SIZE-1:0] key_i;
  logic key_valid_i = 1'b1;
  logic key_ready_o;
  logic [`WORD_SIZE-1:0] hash_o[7:0];
  logic ready_o;
  logic core_ready_o;
  logic done_o;
  
  logic hmac_mode;
  logic [25:0] j = 0;
  logic [511:0]compression;
  logic [63:0] data[130];
  logic [63:0] key[16];
  logic s32;
  string mode, test_str, input_massage;
  typedef enum {test_1,test_2,test_3,test_4,test_5,test_6,test_7} test;
  typedef enum logic[3:0] {sha_256=0,sha_224=1,sha_512=4,sha_384=5,sha_512_256=6,sha_512_224=7,
                HMAC_256=8,HMAC_224=9,HMAC_512=12,HMAC_384=13,HMAC_512_256=14,HMAC_512_224=15} sha_mode;
  test t; sha_mode m; 
    
  lw_hmac uut (
      .opcode_i(opcode_i),
      .clk_i(clk_i), 
      .aresetn_i(aresetn_i), 
      .start_i(start_i),
      .abort_i(abort_i),
      .last_i(last_i),
      .data_valid_i(data_valid_i), 
      .data_i(data_i), 
      .random_i(random_i), 
      .hash_o(hash_o), 
      .ready_o(ready_o),
      .core_ready_o(core_ready_o), 
      .done_o(done_o),
      .key_valid_i(key_valid_i),
      .key_ready_o(key_ready_o),
      .key_i(key_i)
      );
  initial begin
    clk_i = 0;
    forever #5 clk_i = ~clk_i;
  end
  always @(posedge clk_i) random_i <= $random % 4;
  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  task automatic SendBlockData (input [3:0]block_amount);
    int unsigned data_delay = 0, key_delay = 0;
    j = 0;
    while (core_ready_o != 1) @(posedge clk_i);
    if (hmac_mode) begin
      do begin #1;
        start_i = j == 0;
        if (j != 0) opcode_i = 0;
        data_valid_i = j == 0;
        key_valid_i = 1'b1;
        key_i = key[j];
        @(posedge clk_i);
        if (key_valid_i && key_ready_o) j++;
        delay(0, key_delay);
      end while (j < 'd16);
      @(posedge clk_i) begin
        key_valid_i <= 1'b0;
        j = 0;
      end
    end
    
    do begin
      start_i = j == 0 && !hmac_mode;
      if (j != 0) opcode_i = 0;
      data_valid_i = 1'b1;
      data_i = data[j];
      last_i = j == block_amount*16-1;
      @(posedge clk_i);
      if (data_valid_i && ready_o) j++;
      delay(1, data_delay);
    end while (j < block_amount*16);
    @(posedge clk_i) begin #1
      last_i <= 1'b0;
      data_valid_i <= 1'b0;
      j = 0;
    end
    #1 wait (core_ready_o);
    display_output();
    #100;
  endtask
    ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  
  task automatic delay (input logic data, input int unsigned delay);
    repeat(delay) begin #1
      if (data) begin
        data_valid_i = 1'b0;
        data_i = '1;
      end else begin
        key_valid_i = 1'b0;
        key_i = '1;
      end
      start_i = 1'b0;
      last_i = 1'b0;
      @(posedge clk_i);
    end
  endtask
  
  `ifdef CORE_ARCH_S64
  assign hmac_mode = opcode_i[3];
  task automatic display_output();
    if (t==test_1) $display(mode);
    case (m[2:0])
      0: if (hash_o[7:4]==compression[255:0])
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
      1: if (hash_o[7:4]==compression[255:0])
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
       $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
      4: if (hash_o[7:0]==compression)
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
      5: if (hash_o[7:2]==compression[383:0])
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
      6: if (hash_o[7:4]==compression[255:0])
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
      7: if (hash_o[7:4]==compression[255:0])
      $display(test_str, "success!!"); else begin $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);end
    endcase
  endtask
  
  task automatic test_vec_1();
    test_str = "test 1-"; t = test_1;
    input_massage = "NULL";
    data = '{default: 0};
    if (s32) data[0][31] = 1'b1;
    else  data[0][63] = 1'b1;

    if (opcode_i[3]) begin
      data[15] = s32 ? 'd512 : 'd1024;
      case (opcode_i[2:0])
        0: compression = 256'hfd870643c627ffb73a21f861b904e12e1e15ab23d31eaf5ce03dee2f6205a9b0;
        1: compression = 256'ha17c3f1a73654a1fb74c6096d437c17b082d1f6c5b359ed34b6fe1e600000000;
        2: compression = 512'he59cc81631323b25f486646e0b49f58295b3cbd2b8f71389bacc7f8cd6919226452c2bcdb0373005952b2a7c7e5443bf13010e90e0c6ffde49f99804abcd3038;
        3: compression = 384'h9728b939153c6d321b4c3740e21cf14b08c1597186910963898c020a32146709b8c82ed145da6888ce8b1348c74574e7;
        4: compression = 256'heaafb6fc0bd067efe68e2058e0a89337047c148086d523988a538c57b6550e2b;
        5: compression = 256'h4f2fac0ad55f06dfe05e0f9396ab503537bd9cd3a53c91071caca1ee00000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855;
        1: compression = 256'hd14a028c2a3a2bc9476102bb288234c415a2b01f828ea62ac5b3e42f00000000;
        2: compression = 512'hcf83e1357eefb8bdf1542850d66d8007d620e4050b5715dc83f4a921d36ce9ce47d0d13c5d85f2b0ff8318d2877eec2f63b931bd47417a81a538327af927da3e;
        3: compression = 384'h38b060a751ac96384cd9327eb1b1e36a21fdb71114be07434c0cc7bf63f6e1da274edebfe76f65fbd51ad2f14898b95b;
        4: compression = 256'hc672b8d1ef56ed28ab87c3622c5114069bdd3ad7b8f9737498d0c01ecef0967a;
        5: compression = 256'h6ed0dd02806fa89e25de060c19d3ac86cabb87d6a0ddd05c333b84f400000000;
        default: compression = 512'h0;
      endcase
    end
  endtask
  
  task automatic test_vec_2();
    test_str = "test 2-"; t = test_2;
    input_massage = "abc";
    data = '{default: 0};
    data[15] = 64'h0000000000000018;
    data[0] = s32 ? 64'h61626380:64'h6162638000000000;
    if (opcode_i[3]) begin
      data[15] = (s32 ? 'd512:'d1024) + 'h18;
      case (opcode_i[2:0])
        0: compression = 256'h08bc9070da7b1463f1ea0e6993979c5757de84333183a26b69ccc050aed7753e;
        1: compression = 256'h92270d59ae1e0a17d018a2d260c2239b6374dbf581efda635bd35a2500000000;
        2: compression = 512'h62b98f9d34f2ed5b4c286249dd0243a49c43ecda9961235aa775bcbc69c9202edecf1ba36cfab07acc9e4ebb673939b91be567d8f2ac4815765c6f023b034982;
        3: compression = 384'h7e88d1b673a0386b1d17642496312db58d6aa8510e5592646a3e98f7e2de64c3a19aef5901dd50f285e7dca35514d6d3;
        4: compression = 256'h8bd12648ae28b326bc5b25d7d25457b749eafb8d7deee752562b65ce755c8db3;
        5: compression = 256'hfb0b0cb3582a544a33f27fcb9f02d9e60e5b0adaefd70f3a01f29df700000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'hba7816bf8f01cfea414140de5dae2223b00361a396177a9cb410ff61f20015ad;
        1: compression = 256'h23097d223405d8228642a477bda255b32aadbce4bda0b3f7e36c9da700000000;
        2: compression = 512'hddaf35a193617abacc417349ae20413112e6fa4e89a97ea20a9eeee64b55d39a2192992a274fc1a836ba3c23a3feebbd454d4423643ce80e2a9ac94fa54ca49f;
        3: compression = 384'hcb00753f45a35e8bb5a03d699ac65007272c32ab0eded1631a8b605a43ff5bed8086072ba1e7cc2358baeca134c825a7;
        4: compression = 256'h53048e2681941ef99b2e29b76b4c7dabe4c2d0c634fc6d46e0e2f13107e7af23;
        5: compression = 256'h4634270f707b6a54daae7530460842e20e37ed265ceee9a43e8924aa00000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask

  task automatic test_vec_3();
    test_str = "test 3-"; t = test_3;
    if (s32) begin
    input_massage = "abcdbcdecdefdefgefghfghighijhijkijkljklmklmnlmnomnopnopq";
      data = '{default: 0};
      data[31] = 'h1c0;
      data[0:14] = {64'h61626364, 64'h62636465,
                    64'h63646566, 64'h64656667,
                    64'h65666768, 64'h66676869,
                    64'h6768696A, 64'h68696A6B,
                    64'h696A6B6C, 64'h6A6B6C6D,
                    64'h6B6C6D6E, 64'h6C6D6E6F,
                    64'h6D6E6F70, 64'h6E6F7071,
                    64'h80000000};

    end else begin
      input_massage = "abcdefghbcdefghicdefghijdefghijkefghijklfghijklmghijklmnhijklmnoijklmnopjklmnopqklmnopqrlmnopqrsmnopqrstnopqrstu";
      data = '{default: 0};
      data[31] = 'h380;
      data[14][63] = 1'b1;
      data[0:13] = {64'h6162636465666768, 64'h6263646566676869,
                    64'h636465666768696a, 64'h6465666768696a6b,
                    64'h65666768696a6b6c, 64'h666768696a6b6c6d,
                    64'h6768696a6b6c6d6e, 64'h68696a6b6c6d6e6f,
                    64'h696a6b6c6d6e6f70, 64'h6a6b6c6d6e6f7071,
                    64'h6b6c6d6e6f707172, 64'h6c6d6e6f70717273,
                    64'h6d6e6f7071727374, 64'h6e6f707172737475};
    end
    if (opcode_i[3]) begin
      data[31] = s32 ? 'd512 + 'h1c0:'d1024 + 'h380;
      case (opcode_i[2:0])
        0: compression = 256'h615883c8155bcc280a560082d86617444fae38633ccd380b0a24b3314730e841;
        1: compression = 256'hc538385d09aa0ac04abb755b1462b2b3a15dd98f5580d0f97524716a00000000;
        2: compression = 512'h6d9b7df81e01ba42289f0504f538b09d33e97432df6669d7df3c4b5b321bf0fa872303466d020f34aa6852a3a922989a257399be0a7eb52dc074014cfff2090a;
        3: compression = 384'hbd2eb483fbb49d47d5730dbd7d2ea31b426d5f882da2adc8fac5a16ff29a457928dc6b5877cbd636f1a3234089103e6f;
        4: compression = 256'h7324d23123e7d5982d93f338fb0e08ceb7404e88d511d359282664b05b79ab4d;
        5: compression = 256'he0f73d3de8b48ab9225f76b71ddaf632649cf3386af1501a91eda8a600000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'h248d6a61d20638b8e5c026930c3e6039a33ce45964ff2167f6ecedd419db06c1;
        1: compression = 256'h75388b16512776cc5dba5da1fd890150b0c6455cb4f58b195252252500000000;
        2: compression = 512'h8e959b75dae313da8cf4f72814fc143f8f7779c6eb9f7fa17299aeadb6889018501d289e4900f7e4331b99dec4b5433ac7d329eeb6dd26545e96e55b874be909;
        3: compression = 384'h09330c33f71147e83d192fc782cd1b4753111b173b3b05d22fa08086e3b0f712fcc7c71a557e2db966c3e9fa91746039;
        4: compression = 256'h3928e184fb8690f840da3988121d31be65cb9d3ef83ee6146feac861e19b563a;
        5: compression = 256'h23fec5bb94d60b23308192640b0c453335d664734fe40e7268674af900000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask
  
  task automatic test_vec_4();
    test_str = "test 4-"; t = test_4;
    if (s32) input_massage ="rewqiuytsapohgfd;lkjcxz'mbnvf/.,nbedxvium,aw5duinuerfxsbvbastyxmoiuytrewgfdslkjh,mnbvcxzxzaqwsxcedcvrfvbtgbnyhnmujm,rewqiuytsapohgfd;lkjcxz'mbnvf/.,";
    else input_massage = "aaaarewqaaaaiuytaaaasapoaaaahgfdaaaa;lkjaaaacxz'aaaambnvaaaaf/.,aaaanbedaaaaxviuaaaam,awaaaa5duiaaaanueraaaafxsbaaaavbasaaaatyxmaaaaoiuyaaaatrewaaaagfdsaaaalkjhaaaa,mnbaaaavcxzaaaaxzaqaaaawsxcaaaaedcvaaaarfvbaaaatgbnaaaayhnmaaaaujm,aaaarewqaaaaiuytaaaasapoaaaahgfdaaaa;lkjaaaacxz'aaaambnvaaaaf/.,";
    data = '{default: 0};
    data[0:36] = {64'h6161616172657771,    64'h6161616169757974,    64'h616161617361706f,    64'h6161616168676664,
                  64'h616161613b6c6b6a,    64'h6161616163787a27,    64'h616161616d626e76,    64'h61616161662f2e2c,
                  64'h616161616e626564,    64'h6161616178766975,    64'h616161616d2c6177,    64'h6161616135647569,
                  64'h616161616e756572,    64'h6161616166787362,    64'h6161616176626173,    64'h616161617479786d,
                  64'h616161616f697579,    64'h6161616174726577,    64'h6161616167666473,    64'h616161616c6b6a68,
                  64'h616161612c6d6e62,    64'h616161617663787a,    64'h61616161787a6171,    64'h6161616177737863,
                  64'h6161616165646376,    64'h6161616172667662,    64'h616161617467626e,    64'h6161616179686e6d,
                  64'h61616161756a6d2c,    64'h6161616172657771,    64'h6161616169757974,    64'h616161617361706f,
                  64'h6161616168676664,    64'h616161613b6c6b6a,    64'h6161616163787a27,    64'h616161616d626e76,
                  64'h61616161662f2e2c};
      data[47] = s32 ? 64'h4a0 : 64'h940;
      data[37][s32?31:63] = 1'b1;
    if (opcode_i[3]) begin
      data[47] = s32 ? 'd512 + 'h4a0:'d1024 + 'h940;
      case (opcode_i[2:0])
        0: compression = 256'ha80554903afdd812a8b05e110626096e7b647f26df213e80abc596b7f337489a;
        1: compression = 256'hea36672dbce79da3a7308a1992f349920d2db6bfd12abcfe652fc28900000000;
        2: compression = 512'h1de9e6d28842cf76ddb0b73badfcfc9a25d5fafcd743b1f115c0cd271350b0e2043b4e6b8176691d91955166838d54766fce74f9483f2ff15ac5beb9fd8c7606;
        3: compression = 384'hce1b1c442bd3e0985da0b51e307c76d4492a3910d7e5deef9d0b805a444339d1156a44c0c85f42cdd743d0f82a5212c3;
        4: compression = 256'hda976011e6f7c2c17219f8e73025d997ae445d327a281767691ca8a91641c975;
        5: compression = 256'hcd7b4abae8e43a12c788938783eec7b4a53b01b9e44ec1aed375d44300000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'h26d707651fcfe0bcef4e732e3a77a89b312aab802dfdee98fc038036a29283e4;
        1: compression = 256'h0c5cc1d83146f5a32ec721889e9a555476fb506e5627192feeb0143a00000000;
        2: compression = 512'ha8fff1b4852cd61ce420694afea1d19a1e7e217525abd87908713cd38c5488c5f14a9f3a27965db8df4057825c6a859ea72ba587b0cda060c4fda7c5f61cd3e4;
        3: compression = 384'h4b24c0365ffc1119ab358e0d178d5f708bed4a7fd773f81261b48829c77aff9331ea8d6381d3d27abc61941d8d61ffa9;
        4: compression = 256'h6274ebbc8dcf5efee0a597be472eef24097670bf525b9a021ab4e31c225431d9;
        5: compression = 256'h2e34faefa7016ec223c1799f7c01f73de17e8d444828800d6102edc400000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask
  
  task automatic test_vec_5();
    test_str = "test 5-"; t = test_5;
    if (s32) input_massage ="88866d5a04c2b81f579962b7293928a6a2458381ef4f022fc2ec7a72422b275e0f5588e36c63f371a4ddd72d89308a6d1a41e5edced3f805720ecea64f09d21b1059ff90b5b1f5e9ff7f3374da3ded1d47eb9f6562d0bff48974c0234e5be5fa1f571c984c5d4dc8edbd13d4fffc20b5009578b782b7f6b029d1b1b4c7726ef8870d1b9130d967e6b170352e3c1d04579ad3f1207efca01c6d0d4416329e118a66fb0974bac9a026e5511650a4a2a1c10264cf24c38d0c66f3cf3102e2c5be3e69ffd24fcf964f94dcc329543f8be0b67d3ec91547a61ce928ff1e2d1072c1ab9b499dda9a37847747d0011f6457f03dafdce9e23ea6bbbf4371eae2b4278f914ac099c428bdac62d9e0e28a8c97dfd9942a26bb9323b199787ec001a4fc7d8cda3db0928947ddaa9c73dd1a5a496d6e86adaca8ef5b071bda3269f9a31629d8";
    else input_massage = "e6e3f8e688866d5aace56b5104c2b81f2018c313579962b7c6354eca293928a653c3ce94a24583810a4d1749ef4f022fb650afa7c2ec7a727f45199c422b275e0c6676b60f5588e307bd2fe86c63f3712f161f70a4ddd72df9373e2d89308a6df583789d1a41e5edca6ad14eced3f8054d0644ba720ecea679fc057f4f09d21b49e657721059ff90c877faf0b5b1f5e9e0f4e816ff7f3374e41907aada3ded1da34aa42947eb9f651ad3757262d0bff41fca46548974c023a6b97ea34e5be5fa3123ee961f571c98c2163b7f4c5d4dc896c0163dedbd13d403feb51cfffc20b5924ff032009578b71094c54782b7f6b007f9687229d1b1b46fecd110c7726ef8deafb5db870d1b91a3dfecba30d967e624b722a3b170352ea50cb10d3c1d0457ebfc6f9a9ad3f1205daf2cbc7efca01c178bbd696d0d44163e214615329e118ac4f8f82d66fb0974255ec7a0bac9a026bfff2feee5511650aac079fba4a2a1c17c3dafdd0264cf241242500dc38d0c663e56ebc4f3cf31020fdce116e2c5be3ed9d590cb69ffd24f036cb56fcf964f94d4f5c702dcc32954f0dab7533f8be0b6eaae6e6e7d3ec915ec7f4a1347a61ce9af868f7528ff1e2d528add981072c1ab107a9c2f9b499dda34e11d2a9a37847780a2b49647d0011f63e7fd806457f03d5c33fa38afdce9e2fe6f618c3ea6bbbf4e54d9e04371eae2764c1ef7b4278f911027361f4ac099c4fa9d1e0028bdac622b669e27d9e0e28a3d93e0598c97dfd95fa61c62942a26bb2abf21e19323b19923442d99787ec0013f694bf9a4fc7d8cdcdd6339da3db0929af7b8e58947ddaac137331f9c73dd1aa9c62a685a496d6e9991e65286adaca8e9b8263eef5b071bcdaa1882da3269f90cebdb81a31629d8";
    data = '{default: 0};
    data[0:79] = {'he6e3f8e688866d5a, 'hace56b5104c2b81f, 'h2018c313579962b7, 'hc6354eca293928a6,
                  'h53c3ce94a2458381, 'h0a4d1749ef4f022f, 'hb650afa7c2ec7a72, 'h7f45199c422b275e,
                  'h0c6676b60f5588e3, 'h07bd2fe86c63f371, 'h2f161f70a4ddd72d, 'hf9373e2d89308a6d,
                  'hf583789d1a41e5ed, 'hca6ad14eced3f805, 'h4d0644ba720ecea6, 'h79fc057f4f09d21b,
                  'h49e657721059ff90, 'hc877faf0b5b1f5e9, 'he0f4e816ff7f3374, 'he41907aada3ded1d,
                  'ha34aa42947eb9f65, 'h1ad3757262d0bff4, 'h1fca46548974c023, 'ha6b97ea34e5be5fa,
                  'h3123ee961f571c98, 'hc2163b7f4c5d4dc8, 'h96c0163dedbd13d4, 'h03feb51cfffc20b5,
                  'h924ff032009578b7, 'h1094c54782b7f6b0, 'h07f9687229d1b1b4, 'h6fecd110c7726ef8,
                  'hdeafb5db870d1b91, 'ha3dfecba30d967e6, 'h24b722a3b170352e, 'ha50cb10d3c1d0457,
                  'hebfc6f9a9ad3f120, 'h5daf2cbc7efca01c, 'h178bbd696d0d4416, 'h3e214615329e118a,
                  'hc4f8f82d66fb0974, 'h255ec7a0bac9a026, 'hbfff2feee5511650, 'haac079fba4a2a1c1,
                  'h7c3dafdd0264cf24, 'h1242500dc38d0c66, 'h3e56ebc4f3cf3102, 'h0fdce116e2c5be3e,
                  'hd9d590cb69ffd24f, 'h036cb56fcf964f94, 'hd4f5c702dcc32954, 'hf0dab7533f8be0b6,
                  'heaae6e6e7d3ec915, 'hec7f4a1347a61ce9, 'haf868f7528ff1e2d, 'h528add981072c1ab,
                  'h107a9c2f9b499dda, 'h34e11d2a9a378477, 'h80a2b49647d0011f, 'h63e7fd806457f03d,
                  'h5c33fa38afdce9e2, 'hfe6f618c3ea6bbbf, 'h4e54d9e04371eae2, 'h764c1ef7b4278f91,
                  'h1027361f4ac099c4, 'hfa9d1e0028bdac62, 'h2b669e27d9e0e28a, 'h3d93e0598c97dfd9,
                  'h5fa61c62942a26bb, 'h2abf21e19323b199, 'h23442d99787ec001, 'h3f694bf9a4fc7d8c,
                  'hdcdd6339da3db092, 'h9af7b8e58947ddaa, 'hc137331f9c73dd1a, 'ha9c62a685a496d6e,
                  'h9991e65286adaca8, 'he9b8263eef5b071b, 'hcdaa1882da3269f9, 'h0cebdb81a31629d8};
    data[95] = s32 ? 64'ha00 : 64'h1400;
    data[80][s32?31:63] = 1'b1;
    if (opcode_i[3]) begin
      data[95] = s32 ? 'd512 + 'ha00:'d1024 + 'h1400;
      case (opcode_i[2:0])
        0: compression = 256'hda318988b27a1ecda8bc5ccb0f77a5457d8e6221992cb5ff4d7b09dea1b00cbe;
        1: compression = 256'h69efc48a364aebb517f22375bfc5a65a478e39bb881b8c369d9997ee00000000;
        2: compression = 512'h584433b7ee921ca69abb525f5f0f2618d7afe6c561beb67967e23b56e69ad42c6c342eb58e1bf6d0e625c420a57430d5c62dbb48129ebda877e225a76827348c;
        3: compression = 384'he2b957904ccf536ad11a81c3fdd2be197f8a30ae97a951154867be311d330fcedb361821de9aac293a5982d0eb416d19;
        4: compression = 256'ha2630566991fcd58b1d4e28ab048732fcace366b9c566f58de6dec0bb5fa6a6f;
        5: compression = 256'hdf4caa0897f8ffbe256b02a440fabae54a71286c9546ef2f02fdc30c00000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'h826d606f511f043501117d7ae6cf2e797aadeeb86ecd8be7f59335f32ccb0ac3;
        1: compression = 256'h470aea87bd2cb484ee41d38c01693c367c86a8aacb404eacf32130fa00000000;
        2: compression = 512'h172de649b07f51fde7980f0b769d1cc128ab1efb3d8fcd2af603a2becc4f688f5be8a9b600982565d021d5fcf66cdf207e20c3863ba4404b7114636105e2b2fc;
        3: compression = 384'h456109a1ea6b47e0a9289e4eccd3eec9f2e60afe869615816b9a79e86d025809981a1a58ed69ab03c891a4a71fcb85d4;
        4: compression = 256'h4ee2088160129056e0e474ec16993fc572e86eae85f4a4e1f5a105b10efb0181;
        5: compression = 256'h03714a750dacbd8b2c59b257133d6c7d61adc5f6ba647cb365c33f0e00000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask
  
  task automatic test_vec_6();
    test_str = "test 6-"; t= test_6;
    if (s32) input_massage ="d364e8f1545ce324431f92858db5d670dbb90c597149fd94402fbef07d04a3f76e5604c98102eec5adb391582c6758b85ddd03f53b1696b125c71235cf692dd45f260dd4fe1e19759544655511310ce88581166caa512601073ddceaa9a0d3608952ecd51bf2a12ed18ad3d8a246c2098d97d8dc762483c49ce8e1ccb4c7ff8721b765046af02a3b44fa8a4ffb474e3c8dfc121c7a4fcf5cf597b269b8465ed838be2884645a504f251846bd82e8ccdcc7f4296b6995d44fd2b3634322c119a11abdcff594756536f1d217d65dfcc6e48dfe4976865425f17f95f9b420368ea99df22598c33f49b0a9f669485e5661682d698fc973c0e1b4627d53fe417e82be13243d29ef5c950f56cb298cedbffac5899ca76c4e785cf683468eb897aca16e0438df074093b0e177e94d707ebece79fe133407a7f48756c5d112f3de2ff50e";
    else input_massage = "7794cc3dd364e8f1e09d1a01545ce3245507945b431f92855bfc5e6c8db5d6703a70f2a4dbb90c59277e4d9b7149fd943e1f2098402fbef06e91e2bf7d04a3f7d52c59156e5604c9a00c386b8102eec58b4d7516adb391582a2631ae2c6758b8fa14ee1c5ddd03f500deb1fe3b1696b19bdc06a725c71235c19bf174cf692dd4873228985f260dd4df2a943afe1e1975a0376d409544655565e5752911310ce8bbaf26338581166c1ae70046aa512601f6f5cfc0073ddcea1e98d569a9a0d360f1852d1c8952ecd596e6bca81bf2a12e61e26ba9d18ad3d8a25aa131a246c209da976c748d97d8dcddce6ad5762483c463404bdf9ce8e1cc3aa29fe6b4c7ff87e6bf8a6821b76504ba61dea66af02a3b3ff028c444fa8a4f256333e6fb474e3c707b78758dfc121c9f38ecc97a4fcf5c8a0a9995f597b26944a54e5fb8465ed8f327255438be2884e0334b97645a504f42d7fd66251846bd8dfc70da82e8ccdc1ca860d2c7f4296b91353bae6995d44f4a7b69dad2b36343b0fca6e922c119a1ddd0f86d1abdcff5f47084e4947565361394f23af1d217d65342c6285dfcc6e4a39cc4928dfe4976b07d6156865425f1129438387f95f9b44718e6f720368ea9e51cb8289df2259899bb3a2cc33f49b0bde2c64ea9f66948bf9043885e566168a087ce262d698fc99b1eed3273c0e1b4dd477829627d53fe17c16b85417e82bee21ac93e13243d29b9b5cb46ef5c950f420d2c9656cb298c03913407edbffac57db4cbcd899ca76c7b8582b54e785cf692ab7be983468eb82784bbb497aca16e7bfd75590438df07e1c0e7874093b0e1fd73f25d77e94d70f823391d7ebece79f3a929cefe133407aa9cf54fa7f48756712c2ec4c5d112f380077bc3de2ff50e";
    data = '{default: 0};
    data[0:79] = {'h7794cc3dd364e8f1, 'he09d1a01545ce324, 'h5507945b431f9285, 'h5bfc5e6c8db5d670, 
                  'h3a70f2a4dbb90c59, 'h277e4d9b7149fd94, 'h3e1f2098402fbef0, 'h6e91e2bf7d04a3f7, 
                  'hd52c59156e5604c9, 'ha00c386b8102eec5, 'h8b4d7516adb39158, 'h2a2631ae2c6758b8, 
                  'hfa14ee1c5ddd03f5, 'h00deb1fe3b1696b1, 'h9bdc06a725c71235, 'hc19bf174cf692dd4, 
                  'h873228985f260dd4, 'hdf2a943afe1e1975, 'ha0376d4095446555, 'h65e5752911310ce8, 
                  'hbbaf26338581166c, 'h1ae70046aa512601, 'hf6f5cfc0073ddcea, 'h1e98d569a9a0d360, 
                  'hf1852d1c8952ecd5, 'h96e6bca81bf2a12e, 'h61e26ba9d18ad3d8, 'ha25aa131a246c209, 
                  'hda976c748d97d8dc, 'hddce6ad5762483c4, 'h63404bdf9ce8e1cc, 'h3aa29fe6b4c7ff87, 
                  'he6bf8a6821b76504, 'hba61dea66af02a3b, 'h3ff028c444fa8a4f, 'h256333e6fb474e3c, 
                  'h707b78758dfc121c, 'h9f38ecc97a4fcf5c, 'h8a0a9995f597b269, 'h44a54e5fb8465ed8, 
                  'hf327255438be2884, 'he0334b97645a504f, 'h42d7fd66251846bd, 'h8dfc70da82e8ccdc, 
                  'h1ca860d2c7f4296b, 'h91353bae6995d44f, 'h4a7b69dad2b36343, 'hb0fca6e922c119a1, 
                  'hddd0f86d1abdcff5, 'hf47084e494756536, 'h1394f23af1d217d6, 'h5342c6285dfcc6e4, 
                  'ha39cc4928dfe4976, 'hb07d6156865425f1, 'h129438387f95f9b4, 'h4718e6f720368ea9, 
                  'he51cb8289df22598, 'h99bb3a2cc33f49b0, 'hbde2c64ea9f66948, 'hbf9043885e566168, 
                  'ha087ce262d698fc9, 'h9b1eed3273c0e1b4, 'hdd477829627d53fe, 'h17c16b85417e82be, 
                  'he21ac93e13243d29, 'hb9b5cb46ef5c950f, 'h420d2c9656cb298c, 'h03913407edbffac5, 
                  'h7db4cbcd899ca76c, 'h7b8582b54e785cf6, 'h92ab7be983468eb8, 'h2784bbb497aca16e, 
                  'h7bfd75590438df07, 'he1c0e7874093b0e1, 'hfd73f25d77e94d70, 'hf823391d7ebece79, 
                  'hf3a929cefe133407, 'haa9cf54fa7f48756, 'h712c2ec4c5d112f3, 'h80077bc3de2ff50e };
    data[95] = s32 ? 64'ha00 : 64'h1400;
    data[80][s32?31:63] = 1'b1;
                
    if (opcode_i[3]) begin
      data[95] = s32 ? 'd512 + 'ha00:'d1024 + 'h1400;
      case (opcode_i[2:0])
        0: compression = 256'hb418358be947c67ea5056b229cd4f2217042d9c52d37afcae1f95bca1e51a149;
        1: compression = 256'h6927ec1ea452b542606d8ed095ecbc0e83b29e7454b1b0906fd29b1700000000;
        2: compression = 512'ha586e2c3d788d1e56c1354e5bee0154119cc10978a2469d537a36488ff217eb75754a2104b81c7c295a1f89f30563fee343d4a4f76a1c1d99f6a231b7217b5bb;
        3: compression = 384'h2e8901a689d99550b07a2cc075c6ab13278c4ac2665730672c6b48c0ae8eeb2809dbe97ab1a13ec1e5b76124d294548d;
        4: compression = 256'h321b11c590e81bd165ebba578b738132dac992240d4210a9c379bd9e327380d9;
        5: compression = 256'h3e5f8406eba03fc02c05d88553b43216a647831e82a97849c978a39300000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'he23e005624bcc730f352a672e6ddd1500ea787eccd386d71485c7e1c953fb898;
        1: compression = 256'h24468bf42cc037aa0f73c98e717db14c5c01469acfd5dcf49a3b22ca00000000;
        2: compression = 512'h8a953e520970b81d09a8a9d58fc2f27b8f6eb0a487a3ffe4d5cea25be6e15988ffad4ac1e6ade1cd599ee8741a86e80371b0931ce1d0d62ff1ef5586ca579dbd;
        3: compression = 384'h9d4309d012cb1cdc0ed4b58b61cab1700ff7d3cbdba4515d9a9fdfb8592824c8bc9c38ec96957f02082d35eaa98b566c;
        4: compression = 256'h3eee58e304b4013badc17dba36660d9f87333984145cc5b37a4fda4e6bce7ba7;
        5: compression = 256'h75c7b9c42cf08c5c3bd804911f93b9ae1ae615d6998b268beb2cab0200000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask
  
  task automatic test_vec_7();
    test_str = "test 7-"; t= test_7;
    if (s32) input_massage ="010010000111000001011110100110010100010011011010010001001011010011001000000100111000111100110000100000011010000000000001110100101111001010001010110011000001011001110100010101101011001011000111011110110011011001101011110011000001110010000001010001110100010111001100011000010001010011010111011010111100110001000010010000111000000110110101010001010011111011000111100000110011101101111101111010011100001011001111000011111000101000011000010111011110111110001000011110110101011111011010100000101010001011100111010111101001100010111001110101010011010001110010010110011010110011001111100001001011011100011000001101011001000000011100100100110000111001101100100101010100000011111010000001011110101100010111001010001010010011010101010000110010010101110000011011011100100011110001001101011110000101101001010110000110001101101011110010010111111101011010100000111101000010111110111001000101001101010000101011010000001101101011111010011000001011101110101101100010101010011010010101101010110011111000010101011110110111001010001101000010011100101001001111111001100011101100010001011110100111100010011111001000101001111111001101011000000011001100000100001011110010000100001101111010110010010000010011010100110001100001110111000110110000100110011010010011111100010011000000101010000101110001001010001111111000111101001010101001100000100001101110100011111111101110100111000001010100001110001001001111001110110001110110111000100011111100000011111110000000110010011111010011011101101100011110011100011100101101111000000111101101101101101011001000000110110011101101000010111001100000001111111110110010000010100011111100000110001010110000100101010100010111011010111100101111000111010010010100000011111111101101001101100001111111011000111111110100100100000100110000100111011101100000010001010111011000000100101000011010011011010110010101110101101110010011111010111001011100111010000111101010110100000010110000010010000111101111100001110111101100110000000010010011111101001101111011000110000001101101101001110010110100011000101110000110110001001011100100011110010000111100000000111111111011100011011100001110001011110110001101011100010111110000101000111010001100110101100000110101000001111011000001111111111100000100111100111110001110110010000010100110100011011001101100100111111011001111011101111000100011100100110011101101011000101011101100010100101110110001101010111110100110000101011100100001101010010110100010000011010101010011011100010111011111101101101111000110100011000000011001100011111000110010100111100101011011100101110010000011010101111010110011110001111000000111100100101110110010010001001100000111110111100011100010011100011101001000110001011111111000011000010001001111010100001011000011000000011011101100100010010110011101111110000011111001010000010001000011010111001000010111100100101001100110111111010111100010010010001011111011011011100100110101111010010010111011111011100110010110101110010101111101001110111110000000000101010011110111011101011010010010011010000101011100010100101010111011010101110110111100100010111011101000001110000110111110111111001011000101110011111110101011001010010100111111010000011111001001110101011110011101111101000010100110100001101010100000101001001001001000101000101001000110000011010111111110010001111010111110011010011001010001101010100100000010001101101010111010110101000100100111010110100011110001010010000101110000000101110011011101101110110111000110011101110000010000100000001000101110100000000011001110011110000110101100101011110100000010001110010111011000000100110010011110100100000111001101010001000100111110101101111011001011011110001110010000100100010010010110001111000011011101010001101010110110000011000010110001010010000010010111010100011000011001111100100110111110111011001010010111101101110001110100001011100100000000011111000000101010100101100011111001010010010011000110100001110010100001001001100001101100101111010110111100001001010101110001010011110001111101001000110000100001110101111110101101111011111001100101111001101011100";
    else input_massage = "000010101011100001101111111101000100100001110000010111101001100110010100100101011001111101001101010001001101101001000100101101000001001111000000011011000011111011001000000100111000111100110000011101110011010101110000010011011000000110100000000000011101001000111100010011000011000100110101111100101000101011001100000101100100000100111110100101111000110101110100010101101011001011000111110110001110010110100100101001010111101100110110011010111100110000011001110000110101111110110001000111001000000101000111010001010111110101000110000100010010100111001100011000010001010011010111101010000100101010110100011011110110101111001100010000100100001110000101111000001010100110110011100000011011010101000101001111101001100001001110101010010001010011000111100000110011101101111101100100000101011111111110000001111110100111000010110011110000111100011100101111001111001111111101100010100001100001011101111011110000000000000010100010010100000010001000011110110101011111011010011010000111011001101011000111101000001010100010111001110101111001111100011011110010010001001010100110001011100111010101001101001010001101001101001110010000011101110010010110011010110011001111111101101110110111001001000001101000010010110111000110000011010101100011111000011100000000101011100100000001110010010011000011100010101110101000010110111111111101101100100101010100000011111010000110101010110001010001000100000000010111101011000101110010100010000111111100110011010000000100101001001101010101000011001001011101011111100000111001100010000001110000011011011100100011110001110000010000001100001011100100010011010111100001011010010101100000000010000011100011001101100001011000110110101111001001011111111001110001011111010100111101100001011010100000111101000010111110101100100001000011111010100001101110010001010011010100001010110101001000100101000010000011100111000000110110101111101001100000101110010111100011010001011100000011101110101101100010101010011010010110101001100100100101010110000101011010101100111110000101010100100111101101001000111100101000111011011100101000110100001001111100110111000000101011100011111000101001001111111001100011101100111001110011010110100111110100110100010111101001111000100111110010011000100001000011100010100000100010100111111100110101100000001010000000011010101010110011111111001100000100001011110010000100100110110101110001111111000011000011011110101100100100000100110110111110010110000010000111100110010011000110000111011100011011000001000000101101100001011001001100100110011010010011111100010011101100010010000000110000000100000000001010100001011100010010100001101010100010011110010101011101111111100011110100101010100110000110000101000000101101000100101100100001101110100011111111101110000011010111000100100111111101001001110000010101000011100010010010110101101011001010110100110001010011110011101100011101101110000111110111111011110110110110011110001111110000001111111000000011111110110111010001110010000001100010011111010011011101101100011110111011010100111111100111000000100111000111001011011110000001111010111001001101100110011110110010110110110110101100100000011011111001110101110010110001011110110011101101000010111001100000001110001111101110101111010001111101111111101100100000101000111111001101010111011011101010011101001000011000101011000010010101010001000010011111110101001001000101110111011010111100101111000111010000001011110010001011001110111101100101000000111111111011010011011011000101001110111111011000111010000111111101100011111111010010111001101110110000111101100010000100000100110000100111011101100010010001100100110100011100110011000100010101110110000001001010000010111011110111010110011100001001101001101101011001010111010110110111011100010111000010100100001110010011111010111001011100111010111111011000101100100101100110100001111010101101000000101100000100010010100101010011101111001001001000011110111110000111011110011011011100010110101111000000101100110000000010010011111101001111001110100100010010011011000001011101011011000110000001101101100011011011110001001111101011010010011100000010110100011000101110111100000110101110010111011001100001101100010010111001000111100101110010100100100101100111000000000011110000000011111111101110001100101010011101001111110011100111011100001110001011110110001101000110101011010000100001010111000111000101111100001010001110100010011001110001101000010010101001110011010110000011010100000111101001001001111011101111100010110011000001111111111100000100111100101100000110101101011011010101011111100011101100100000101001101001111000100011011100000000000011001101100110110010011111101100110001011111110010000011101110001011011101111000100011100100110011010111101011001101001001111101111011010110001010111011000101001010110010100010111010011110010100111011000110101011111010011000011010010110101001000111100011011101011100100001101010010110100010101110111011110011110100011100110000110101010100110111000101110101100001010101100011111001011000111110110110111100011010001100001100110000011001001111111100100100011001100011111000110010100111000000011001100111101110000000011001010110111001011100100000110101110010111110100000010011011011010111101011001111000111100000011011110000001011010111111011001011100100101110110010010001001100011001100011011000010111001010000001111101111000111000100111000111010000011000110000001000000111110100100011000101111111100001101010100110111001100110101001110000010001001111010100001011000011111100001111001010000111111000000000000110111011001000100101100110000111110011011101101100011100110111111000001111100101000001000000100111111100111100001000011101000011010111001000010111100100011010001100000101000101000010011010011001101111110101111000100110100000111001011111001110100011001000101111101101101110010011011011100011111110110011011110101101111010010010111011111011100110101000000100010000111100000111010101101011100101011111010011101111000001110111001111101010100111111000000000010101001111011101110110011001010101000101010101001001011010010010011010000101011100000010101001000001001111111100010101001010101110110101011101101111000000111100000111100110011010110010001011101110100000111000010010101111110111000000110100100110111110111111001011000101110011001011101010001111010010000100001111101010110010100101001111110110000000101110001110010101110011000001111100100111010101111001110001011011000001000100010110010101111101000010100110100001101010111011101100101111011100101001011000001010010010010010001010001001110000000111000011001100101111100100011000001101011111111001001111001011111001110000011100000101111010111110011010011001010001111001001000010100111001010001011010101001000000100011011010101111010110011101110100001111000110101011010100010010011101011010001011110011001011011111101011000111110001010010000101110000000101011000101110010001001100001101101100110111011011011100011001110101000111000110010011111111101110110000010000100000001000101110101010011100001100111011000001111100000000110011100111100001101011010010101001010011010000011100010010101111010000001000111001011111010111111100011100111011011011011000000100110010011110100100001011000100101010000111100001101001110011010100010001001111101011110011100010100001101100100100110111101100101101111000111001000001110101001111010100101111011100100100010010010110001111000011011100001010001011100101011100011011010100011010101101100000110000000110110111111110010001001100011011000101001000001001011101010001000101011100110000011010100101011000011001111100100110111110110110111101000110100011010111000110110010100101111011011100011101101111001000110000110111101101000000101110010000000001111100000010110100100100101101000001111001101010100101100011111001010010011001110001100010101011110101100100110001101000011100101000010010010101010110001101100110010010010110000110110010111101011011110010001100111011001000001100001111001001010101110001010011110001110010010110100000001010000001010011010010001100001000011101011111011101011100111101111101101101011010110111101111100110010111100111111010010100110000000001000011101011100";
    data[0:126] = { 'h0ab86ff448705e99, 'h94959f4d44da44b4, 'h13c06c3ec8138f30, 'h7735704d81a001d2, 
                    'h3c4c3135f28acc16, 'h413e978d7456b2c7, 'hd8e5a4a57b366bcc, 'h19c35fb11c814745, 
                    'h7d461129cc6114d7, 'ha84ab46f6bcc4243, 'h85e0a9b381b5453e, 'h984ea914c7833b7d, 
                    'h9057fe07e9c2cf0f, 'h1cbcf3fd8a185def, 'h00028940887b57da, 'h68766b1e82a2e75e, 
                    'h7c6f244a98b9d534, 'ha34d39077259accf, 'hf6edc90684b71835, 'h63e1c02b901c930e, 
                    'h2ba85bff6c9540fa, 'h1aac511005eb1728, 'h87f33404a4d54325, 'hd7e0e620706dc8f1, 
                    'hc1030b9135e16958, 'h020e3361636bc97f, 'h9c5f53d85a83d0be, 'hb210fa86e45350ad, 
                    'h489420e7036be982, 'he5e345c0eeb62a9a, 'h5a99255856acf855, 'h27b48f28edca3427, 
                    'hcdc0ae3e293f98ec, 'he735a7d345e9e27c, 'h988438a08a7f3580, 'ha01aab3fcc10bc84, 
                    'h9b5c7f0c37ac904d, 'hbe5821e64c61dc6c, 'h102d859326693f13, 'hb120301002a17128, 
                    'h6a89e55dfe3d2a98, 'h6140b44b21ba3fee, 'h0d7127f49c150e24, 'hb5acad314f3b1db8, 
                    'h7dfbdb678fc0fe03, 'hfb74720627d376c7, 'hbb53f9c09c72de07, 'hae4d99ecb6dac81b, 
                    'he75cb17b3b42e603, 'h8fbaf47dfec828fc, 'hd5dba9d218ac2551, 'h09fd491776bcbc74, 
                    'h0bc8b3bd940ffb4d, 'hb14efd8e87f63fd2, 'he6ec3d8841309dd8, 'h91934733115d8128, 
                    'h2ef759c269b595d6, 'hddc5c290e4fae5ce, 'hbf62c96687ab40b0, 'h44a54ef2487be1de, 
                    'h6dc5af02cc024fd3, 'hce9126c175b181b6, 'h36f13eb49c0b462e, 'hf06b97661b12e479, 
                    'h729259c00f00ffb8, 'hca9d3f39dc38bd8d, 'h1ab4215c717c28e8, 'h99c684a9cd60d41e, 
                    'h927bbe2cc1ffc13c, 'hb06b5b55f8ec829a, 'h788dc003366c9fb3, 'h17f20ee2dde23933, 
                    'h5eb349f7b58aec52, 'hb28ba794ec6afa61, 'ha5a91e375c86a5a2, 'hbbbcf4730d54dc5d, 
                    'h61563e58fb6f1a30, 'hcc193fc9198f8ca7, 'h0199ee0195b9720d, 'h72fa04db5eb3c781, 
                    'hbc0b5fb2e4bb244c, 'h663617281f78e271, 'hd0630207d2317f86, 'ha9b99a9c113d42c3, 
                    'hf0f287e001bb2259, 'h87cddb1cdf83e504, 'h09fcf087435c85e4, 'h68c14509a66fd789, 
                    'ha0e5f3a322fb6e4d, 'hb8fecdeb7a4bbee6, 'ha0443c1d5ae57d3b, 'hc1dcfaa7e0054f77, 
                    'h665515525a49a15c, 'h0a904ff152aed5db, 'hc0f0799ac8bba0e1, 'h2bf70349befcb173, 
                    'h2ea3d210fab294fd, 'h80b8e57307c9d5e7, 'h16c111657d0a686a, 'heecbdca5829248a2, 
                    'h701c332f91835fe4, 'hf2f9c1c17af9a651, 'he4853945aa408dab, 'hd67743c6ad449d68, 
                    'hbccb7eb1f1485c05, 'h62e44c36cddb719d, 'h47193feec10808ba, 'ha70cec1f00ce786b, 
                    'h4a94d0712bd02397, 'hd7f1cedb604c9e90, 'hb12a1e1a735113eb, 'hce286c937b2de390, 
                    'h753d4bdc91258f0d, 'hc28b95c6d46ad830, 'h1b7f9131b14825d4, 'h457306a5619f26fb, 
                    'h6f468d71b297b71d, 'hbc8c37b40b9007c0, 'hb492d079aa58f949, 'h9c62af5931a1ca12, 
                    'h5563664961b2f5bc, 'h8cec830f255c53c7, 'h25a02814d230875f, 'h75cf7db5adef9979, 
                    'hfa530043ae400000, 'h0000000000000000, 'h0000000000000000 };
                    
    data[127] = s32 ? 64'hf89 : 64'h1f29;
    if (opcode_i[3]) begin
    data[127] = s32 ? 'd512 + 'hf89:'d1024 + 'h1f29;
      case (opcode_i[2:0])
        0: compression = 256'h4820a4a4c044b523a5c292556b0d89125df0a0a6da59a78b953571bf58d6d884;
        1: compression = 256'h44d0c31c0db1388e9c23c4859e239824bdf29059c5a812c3ea501f3900000000;
        2: compression = 512'h068e5203823a9fdd4e7a4d4ec477b0f496ac3b68ecbca43f959aeb12f358bf8c714a1e56f485b73552a0fe339d34f8095c8b2d03c5f5549dfcfc13c78cefaead;
        3: compression = 384'hb7a19e9a88813c13216d96e8a728ab2982051658a54aa333af256a032fe3ad647ad7c328aa793d34087269e845aed5d6;
        4: compression = 256'hf01c2ff12e385cf145c639de06b6035c3c3085669df18f753eb03c0f2ccc9cde;
        5: compression = 256'h30c4e5e1100ad299231eeb7a5a81dfb56ac2e335223fe00e24678c9d00000000;
        default: compression = 512'h0;
      endcase
    end else begin
      case (opcode_i[2:0])
        0: compression = 256'h0637697e16c69aaf54c92a0a4338ba4318235f7ca65937afaf39e5387e06784b;
        1: compression = 256'hb1d2c4905656d571f7ef0806f590be218c814f386ab117310a8d381800000000;
        2: compression = 512'hae756d6fbe7568d68a1ec8fa14c3e101d3dc792befb727545b6001c0969dbf0eb14a1c4f5ece012d17204ad8eb4c440ca4692efb41752e015c3a6d2e7459503f;
        3: compression = 384'hd20d1900403e6e43b00ecd1aa32b1828ed17444d26bb1b7fbfdcc8b98660f7f50ea761e5a3f110c8b2f4d88805466427;
        4: compression = 256'he3ac5bd18a330626b9c0c61961897f4b930e331f3b3ac7ac7cbd1c9fec22735a;
        5: compression = 256'h2c773e64026a633934a35466a2e3db0e7e4e2b5eb2330468a0815c9600000000;
        default: compression = 512'h0;
      endcase
    end
  #1; endtask
  task automatic assigning_key();
    key[0:15] = { 64'h07f089fd09a09c09, 64'h890b9089c989a090,
                  64'h4542345f23b432e2, 64'ha98b09c98000323f,
                  64'h089b977987c79a90, 64'hb4c6ba9908f0ff32,
                  64'h665253463225656e, 64'h62546a453326234f,
                  64'h9809b908ca889df0, 64'h6877a9d980bc09a3,
                  64'h43525245bc54d2af, 64'h6c2345d34b23c26e,
                  64'h624352e332bb2af4, 64'h4525232f23e2a24c,
                  64'h253456324f5233c5, 64'ha9877b9899c7689e };
  #1; endtask
  
  task automatic assigning_simple_key();
    key[0:15] = { 64'hc, 64'hd,
                  64'ha, 64'hb,
                  64'h8, 64'h9,
                  64'h90, 64'h80,
                  64'hf0, 64'he0,
                  64'hd0, 64'hc0,
                  64'hc00, 64'hd00,
                  64'ha00, 64'hb0f };
  #1; endtask
  task automatic reseting();
    aresetn_i <= 0; #20
    aresetn_i <= 1;
  endtask
  
  assign s32 = opcode_i[2:1]==2'b00;
 
  task automatic assigning_title();#1
    case (opcode_i)
      0: begin mode = "sha 256: "; m = sha_256; end
      1: begin mode = "sha 244: "; m = sha_224; end
      2: begin mode = "sha 512: "; m = sha_512; end
      3: begin mode = "sha 384: "; m = sha_384; end
      4: begin mode = "sha 512/256: "; m = sha_512_256; end
      5: begin mode = "sha 512/244: "; m = sha_512_224; end
      8: begin mode = "HMAC 256: "; m = HMAC_256; end
      9: begin mode = "HMAC 244: "; m = HMAC_224; end
      10: begin mode = "HMAC 512: "; m = HMAC_512; end
      11: begin mode = "HMAC 384: "; m = HMAC_384; end
      12: begin mode = "HMAC 512/256: "; m = HMAC_512_256; end
      13: begin mode = "HMAC 512/244: "; m = HMAC_512_224; end
    endcase
  endtask

  task automatic running_tests(input [3:0] opcode);
    #1opcode_i = opcode; assigning_title(); test_vec_1(); SendBlockData(1); // 1 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_2(); SendBlockData(1); // 1 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_3(); SendBlockData(2); // 2 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_4(); SendBlockData(3); // 3 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_5(); SendBlockData(6); // 5 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_6(); SendBlockData(6); // 6 Block data
    #1opcode_i = opcode; assigning_title(); test_vec_7(); SendBlockData(8); // 8 Block data
    $display();
    if (mode == "sha 512/244: ") begin
      $display("/////////////////////////////////////////////////////////");
      $display();
    end
  endtask

  //////////////////////////////////////////////////////
  initial begin
    reseting();
    ////////////////////////////////////////////////////
//    assigning_simple_key();
    assigning_key();
    
    running_tests(0);//SHA-256
    running_tests(1);//SHA-224
    running_tests(2);//SHA-512
    running_tests(3);//SHA-384
    running_tests(4);//SHA-512/256
    running_tests(5);//SHA-512/224
    reseting();
    running_tests(8);//HMAC-256
    running_tests(9);//HMAC-224
    running_tests(10);//HMAC-512
    running_tests(11);//HMAC-384
    running_tests(12);//HMAC-512/256
    running_tests(13);//HMAC-512/224
  end
    ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 
 `else `ifdef CORE_ARCH_S32 
 
  assign hmac_mode = opcode_i[1];
  task automatic display_output();
    if (t==test_1) $display(mode);
    if (hash_o[7:0]==compression) begin
      $display(test_str, "success!!");
    end else begin
      $display(test_str, "failed :(  massage input is:");
      $display(input_massage); $display("The output is: %h", hash_o[7:0]);
    end
  endtask
  
  task automatic test_vec_1();
    test_str = "test 1-"; t = test_1;
    input_massage = "NULL";
    data[0:15] = {32'h80000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000,
                  32'h00000000, 32'h00000000};
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'ha17c3f1a73654a1fb74c6096d437c17b082d1f6c5b359ed34b6fe1e600000000:
        256'hfd870643c627ffb73a21f861b904e12e1e15ab23d31eaf5ce03dee2f6205a9b0;
        data[15] = 'd512;
    end else begin
        compression = opcode_i[0] ?
        256'hd14a028c2a3a2bc9476102bb288234c415a2b01f828ea62ac5b3e42f00000000:
        256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855;
    end
  endtask
  
  task automatic test_vec_2();
  test_str = "test 2-"; t = test_2;
  input_massage = "abc";
      data[0:15] = {32'h61626380, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000000,
                    32'h00000000, 32'h00000018};
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'h92270d59ae1e0a17d018a2d260c2239b6374dbf581efda635bd35a2500000000:
        256'h08bc9070da7b1463f1ea0e6993979c5757de84333183a26b69ccc050aed7753e;
        data[15] = 'd512 + 'h18;
    end else begin
        compression = opcode_i[0] ?
        256'h23097d223405d8228642a477bda255b32aadbce4bda0b3f7e36c9da700000000:
        256'hba7816bf8f01cfea414140de5dae2223b00361a396177a9cb410ff61f20015ad;
    end
  #1; endtask

  task automatic test_vec_3();
  test_str = "test 3-"; t = test_3;
    input_massage = "abcdbcdecdefdefgefghfghighijhijkijkljklmklmnlmnomnopnopq";
      data[0:31] = {'h61626364, 'h62636465,
                    'h63646566, 'h64656667,
                    'h65666768, 'h66676869,
                    'h6768696A, 'h68696A6B,
                    'h696A6B6C, 'h6A6B6C6D,
                    'h6B6C6D6E, 'h6C6D6E6F,
                    'h6D6E6F70, 'h6E6F7071,
                    'h80000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h00000000,
                    'h00000000, 'h000001c0 };
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'hc538385d09aa0ac04abb755b1462b2b3a15dd98f5580d0f97524716a00000000:
        256'h615883c8155bcc280a560082d86617444fae38633ccd380b0a24b3314730e841;
    data[31] = 'd512 + 'h1c0;
    end else begin
        compression = opcode_i[0] ?
        256'h75388b16512776cc5dba5da1fd890150b0c6455cb4f58b195252252500000000:
        256'h248d6a61d20638b8e5c026930c3e6039a33ce45964ff2167f6ecedd419db06c1;
    end
  #1; endtask
  
  task automatic test_vec_4();
  test_str = "test 4-"; t = test_4;
  input_massage ="rewqiuytsapohgfd;lkjcxz'mbnvf/.,nbedxvium,aw5duinuerfxsbvbastyxmoiuytrewgfdslkjh,mnbvcxzxzaqwsxcedcvrfvbtgbnyhnmujm,rewqiuytsapohgfd;lkjcxz'mbnvf/.,";
    data[0:47] = {'h72657771,    'h69757974,    'h7361706f,    'h68676664,
                  'h3b6c6b6a,    'h63787a27,    'h6d626e76,    'h662f2e2c,
                  'h6e626564,    'h78766975,    'h6d2c6177,    'h35647569,
                  'h6e756572,    'h66787362,    'h76626173,    'h7479786d,
                  'h6f697579,    'h74726577,    'h67666473,    'h6c6b6a68,
                  'h2c6d6e62,    'h7663787a,    'h787a6171,    'h77737863,
                  'h65646376,    'h72667662,    'h7467626e,    'h79686e6d,
                  'h756a6d2c,    'h72657771,    'h69757974,    'h7361706f,
                  'h68676664,    'h3b6c6b6a,    'h63787a27,    'h6d626e76,
                  'h662f2e2c,    'h80000000,    'h00000000,    'h00000000,
                  'h00000000,    'h00000000,    'h00000000,    'h00000000,
                  'h00000000,    'h00000000,    'h00000000,    'h000004a0  };
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'hea36672dbce79da3a7308a1992f349920d2db6bfd12abcfe652fc28900000000:
        256'ha80554903afdd812a8b05e110626096e7b647f26df213e80abc596b7f337489a;
        data[47] = 'd512 + 'h4a0;
    end else begin
        compression = opcode_i[0] ?
        256'h0c5cc1d83146f5a32ec721889e9a555476fb506e5627192feeb0143a00000000:
        256'h26d707651fcfe0bcef4e732e3a77a89b312aab802dfdee98fc038036a29283e4;
    end
  #1; endtask
  
  task automatic test_vec_5();
  test_str = "test 5-"; t = test_5;
    input_massage ="88866d5a04c2b81f579962b7293928a6a2458381ef4f022fc2ec7a72422b275e0f5588e36c63f371a4ddd72d89308a6d1a41e5edced3f805720ecea64f09d21b1059ff90b5b1f5e9ff7f3374da3ded1d47eb9f6562d0bff48974c0234e5be5fa1f571c984c5d4dc8edbd13d4fffc20b5009578b782b7f6b029d1b1b4c7726ef8870d1b9130d967e6b170352e3c1d04579ad3f1207efca01c6d0d4416329e118a66fb0974bac9a026e5511650a4a2a1c10264cf24c38d0c66f3cf3102e2c5be3e69ffd24fcf964f94dcc329543f8be0b67d3ec91547a61ce928ff1e2d1072c1ab9b499dda9a37847747d0011f6457f03dafdce9e23ea6bbbf4371eae2b4278f914ac099c428bdac62d9e0e28a8c97dfd9942a26bb9323b199787ec001a4fc7d8cda3db0928947ddaa9c73dd1a5a496d6e86adaca8ef5b071bda3269f9a31629d8";
  data[0:95] = {'h88866d5a, 'h04c2b81f, 'h579962b7, 'h293928a6,
                'ha2458381, 'hef4f022f, 'hc2ec7a72, 'h422b275e,
                'h0f5588e3, 'h6c63f371, 'ha4ddd72d, 'h89308a6d,
                'h1a41e5ed, 'hced3f805, 'h720ecea6, 'h4f09d21b,
                'h1059ff90, 'hb5b1f5e9, 'hff7f3374, 'hda3ded1d,
                'h47eb9f65, 'h62d0bff4, 'h8974c023, 'h4e5be5fa,
                'h1f571c98, 'h4c5d4dc8, 'hedbd13d4, 'hfffc20b5,
                'h009578b7, 'h82b7f6b0, 'h29d1b1b4, 'hc7726ef8,
                'h870d1b91, 'h30d967e6, 'hb170352e, 'h3c1d0457,
                'h9ad3f120, 'h7efca01c, 'h6d0d4416, 'h329e118a,
                'h66fb0974, 'hbac9a026, 'he5511650, 'ha4a2a1c1,
                'h0264cf24, 'hc38d0c66, 'hf3cf3102, 'he2c5be3e,
                'h69ffd24f, 'hcf964f94, 'hdcc32954, 'h3f8be0b6,
                'h7d3ec915, 'h47a61ce9, 'h28ff1e2d, 'h1072c1ab,
                'h9b499dda, 'h9a378477, 'h47d0011f, 'h6457f03d,
                'hafdce9e2, 'h3ea6bbbf, 'h4371eae2, 'hb4278f91,
                'h4ac099c4, 'h28bdac62, 'hd9e0e28a, 'h8c97dfd9,
                'h942a26bb, 'h9323b199, 'h787ec001, 'ha4fc7d8c,
                'hda3db092, 'h8947ddaa, 'h9c73dd1a, 'h5a496d6e,
                'h86adaca8, 'hef5b071b, 'hda3269f9, 'ha31629d8,
                
                'h80000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000a00 };
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'h69efc48a364aebb517f22375bfc5a65a478e39bb881b8c369d9997ee00000000:
        256'hda318988b27a1ecda8bc5ccb0f77a5457d8e6221992cb5ff4d7b09dea1b00cbe;
        data[95] = 'd512 + 'ha00;
    end else begin
        compression = opcode_i[0] ?
        256'h470aea87bd2cb484ee41d38c01693c367c86a8aacb404eacf32130fa00000000:
        256'h826d606f511f043501117d7ae6cf2e797aadeeb86ecd8be7f59335f32ccb0ac3;
    end
  #1; endtask
  
  task automatic test_vec_6();
  test_str = "test 6-"; t= test_6;
    input_massage ="d364e8f1545ce324431f92858db5d670dbb90c597149fd94402fbef07d04a3f76e5604c98102eec5adb391582c6758b85ddd03f53b1696b125c71235cf692dd45f260dd4fe1e19759544655511310ce88581166caa512601073ddceaa9a0d3608952ecd51bf2a12ed18ad3d8a246c2098d97d8dc762483c49ce8e1ccb4c7ff8721b765046af02a3b44fa8a4ffb474e3c8dfc121c7a4fcf5cf597b269b8465ed838be2884645a504f251846bd82e8ccdcc7f4296b6995d44fd2b3634322c119a11abdcff594756536f1d217d65dfcc6e48dfe4976865425f17f95f9b420368ea99df22598c33f49b0a9f669485e5661682d698fc973c0e1b4627d53fe417e82be13243d29ef5c950f56cb298cedbffac5899ca76c4e785cf683468eb897aca16e0438df074093b0e177e94d707ebece79fe133407a7f48756c5d112f3de2ff50e";
  data[0:95] = {'hd364e8f1, 'h545ce324, 'h431f9285, 'h8db5d670,
                'hdbb90c59, 'h7149fd94, 'h402fbef0, 'h7d04a3f7,
                'h6e5604c9, 'h8102eec5, 'hadb39158, 'h2c6758b8,
                'h5ddd03f5, 'h3b1696b1, 'h25c71235, 'hcf692dd4,
                'h5f260dd4, 'hfe1e1975, 'h95446555, 'h11310ce8,
                'h8581166c, 'haa512601, 'h073ddcea, 'ha9a0d360,
                'h8952ecd5, 'h1bf2a12e, 'hd18ad3d8, 'ha246c209,
                'h8d97d8dc, 'h762483c4, 'h9ce8e1cc, 'hb4c7ff87,
                'h21b76504, 'h6af02a3b, 'h44fa8a4f, 'hfb474e3c,
                'h8dfc121c, 'h7a4fcf5c, 'hf597b269, 'hb8465ed8,
                'h38be2884, 'h645a504f, 'h251846bd, 'h82e8ccdc,
                'hc7f4296b, 'h6995d44f, 'hd2b36343, 'h22c119a1,
                'h1abdcff5, 'h94756536, 'hf1d217d6, 'h5dfcc6e4,
                'h8dfe4976, 'h865425f1, 'h7f95f9b4, 'h20368ea9,
                'h9df22598, 'hc33f49b0, 'ha9f66948, 'h5e566168,
                'h2d698fc9, 'h73c0e1b4, 'h627d53fe, 'h417e82be,
                'h13243d29, 'hef5c950f, 'h56cb298c, 'hedbffac5,
                'h899ca76c, 'h4e785cf6, 'h83468eb8, 'h97aca16e,
                'h0438df07, 'h4093b0e1, 'h77e94d70, 'h7ebece79,
                'hfe133407, 'ha7f48756, 'hc5d112f3, 'hde2ff50e,
                                
                'h80000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000000,
                'h00000000, 'h00000000, 'h00000000, 'h00000a00 };
                
    if (opcode_i[1]) begin
        compression = opcode_i[0] ?
        256'h6927ec1ea452b542606d8ed095ecbc0e83b29e7454b1b0906fd29b1700000000:
        256'hb418358be947c67ea5056b229cd4f2217042d9c52d37afcae1f95bca1e51a149;
        data[95] = 'd512 + 'ha00;
    end else begin
        compression = opcode_i[0] ?
        256'h24468bf42cc037aa0f73c98e717db14c5c01469acfd5dcf49a3b22ca00000000:
        256'he23e005624bcc730f352a672e6ddd1500ea787eccd386d71485c7e1c953fb898;
    end
  #1; endtask
  
  task automatic test_vec_7();
  test_str = "test 7-"; t= test_7;
    input_massage ="010010000111000001011110100110010100010011011010010001001011010011001000000100111000111100110000100000011010000000000001110100101111001010001010110011000001011001110100010101101011001011000111011110110011011001101011110011000001110010000001010001110100010111001100011000010001010011010111011010111100110001000010010000111000000110110101010001010011111011000111100000110011101101111101111010011100001011001111000011111000101000011000010111011110111110001000011110110101011111011010100000101010001011100111010111101001100010111001110101010011010001110010010110011010110011001111100001001011011100011000001101011001000000011100100100110000111001101100100101010100000011111010000001011110101100010111001010001010010011010101010000110010010101110000011011011100100011110001001101011110000101101001010110000110001101101011110010010111111101011010100000111101000010111110111001000101001101010000101011010000001101101011111010011000001011101110101101100010101010011010010101101010110011111000010101011110110111001010001101000010011100101001001111111001100011101100010001011110100111100010011111001000101001111111001101011000000011001100000100001011110010000100001101111010110010010000010011010100110001100001110111000110110000100110011010010011111100010011000000101010000101110001001010001111111000111101001010101001100000100001101110100011111111101110100111000001010100001110001001001111001110110001110110111000100011111100000011111110000000110010011111010011011101101100011110011100011100101101111000000111101101101101101011001000000110110011101101000010111001100000001111111110110010000010100011111100000110001010110000100101010100010111011010111100101111000111010010010100000011111111101101001101100001111111011000111111110100100100000100110000100111011101100000010001010111011000000100101000011010011011010110010101110101101110010011111010111001011100111010000111101010110100000010110000010010000111101111100001110111101100110000000010010011111101001101111011000110000001101101101001110010110100011000101110000110110001001011100100011110010000111100000000111111111011100011011100001110001011110110001101011100010111110000101000111010001100110101100000110101000001111011000001111111111100000100111100111110001110110010000010100110100011011001101100100111111011001111011101111000100011100100110011101101011000101011101100010100101110110001101010111110100110000101011100100001101010010110100010000011010101010011011100010111011111101101101111000110100011000000011001100011111000110010100111100101011011100101110010000011010101111010110011110001111000000111100100101110110010010001001100000111110111100011100010011100011101001000110001011111111000011000010001001111010100001011000011000000011011101100100010010110011101111110000011111001010000010001000011010111001000010111100100101001100110111111010111100010010010001011111011011011100100110101111010010010111011111011100110010110101110010101111101001110111110000000000101010011110111011101011010010010011010000101011100010100101010111011010101110110111100100010111011101000001110000110111110111111001011000101110011111110101011001010010100111111010000011111001001110101011110011101111101000010100110100001101010100000101001001001001000101000101001000110000011010111111110010001111010111110011010011001010001101010100100000010001101101010111010110101000100100111010110100011110001010010000101110000000101110011011101101110110111000110011101110000010000100000001000101110100000000011001110011110000110101100101011110100000010001110010111011000000100110010011110100100000111001101010001000100111110101101111011001011011110001110010000100100010010010110001111000011011101010001101010110110000011000010110001010010000010010111010100011000011001111100100110111110111011001010010111101101110001110100001011100100000000011111000000101010100101100011111001010010010011000110100001110010100001001001100001101100101111010110111100001001010101110001010011110001111101001000110000100001110101111110101101111011111001100101111001101011100";
    data[0:127] = {'h48705e99, 'h44da44b4, 'hc8138f30, 'h81a001d2, 'hf28acc16, 'h7456b2c7,
                   'h7b366bcc, 'h1c814745, 'hcc6114d7, 'h6bcc4243, 'h81b5453e, 'hc7833b7d,
                   'he9c2cf0f, 'h8a185def, 'h887b57da, 'h82a2e75e, 'h98b9d534, 'h7259accf,
                   'h84b71835, 'h901c930e, 'h6c9540fa, 'h05eb1728, 'ha4d54325, 'h706dc8f1,
                   'h35e16958, 'h636bc97f, 'h5a83d0be, 'he45350ad, 'h036be982, 'heeb62a9a,
                   'h56acf855, 'hedca3427, 'h293f98ec, 'h45e9e27c, 'h8a7f3580, 'hcc10bc84,
                   'h37ac904d, 'h4c61dc6c, 'h26693f13, 'h02a17128, 'hfe3d2a98, 'h21ba3fee,
                   'h9c150e24, 'h4f3b1db8, 'h8fc0fe03, 'h27d376c7, 'h9c72de07, 'hb6dac81b,
                   'h3b42e603, 'hfec828fc, 'h18ac2551, 'h76bcbc74, 'h940ffb4d, 'h87f63fd2,
                   'h41309dd8, 'h115d8128, 'h69b595d6, 'he4fae5ce, 'h87ab40b0, 'h487be1de,
                   'hcc024fd3, 'h75b181b6, 'h9c0b462e, 'h1b12e479, 'h0f00ffb8, 'hdc38bd8d,
                   'h717c28e8, 'hcd60d41e, 'hc1ffc13c, 'hf8ec829a, 'h366c9fb3, 'hdde23933,
                   'hb58aec52, 'hec6afa61, 'h5c86a5a2, 'h0d54dc5d, 'hfb6f1a30, 'h198f8ca7,
                   'h95b9720d, 'h5eb3c781, 'he4bb244c, 'h1f78e271, 'hd2317f86, 'h113d42c3,
                   'h01bb2259, 'hdf83e504, 'h435c85e4, 'ha66fd789, 'h22fb6e4d, 'h7a4bbee6,
                   'h5ae57d3b, 'he0054f77, 'h5a49a15c, 'h52aed5db, 'hc8bba0e1, 'hbefcb173,
                   'hfab294fd, 'h07c9d5e7, 'h7d0a686a, 'h829248a2, 'h91835fe4, 'h7af9a651,
                   'haa408dab, 'had449d68, 'hf1485c05, 'hcddb719d, 'hc10808ba, 'h00ce786b,
                   'h2bd02397, 'h604c9e90, 'h735113eb, 'h7b2de390, 'h91258f0d, 'hd46ad830,
                   'hb14825d4, 'h619f26fb, 'hb297b71d, 'h0b9007c0, 'haa58f949, 'h31a1ca12,
                   'h61b2f5bc, 'h255c53c7, 'hd230875f, 'hadef9979, 'hae400000, 'h00000000,
                   'h00000000, 'h00000f89 };
    if (opcode_i[1]) begin
      compression = opcode_i[0] ?
      256'h44d0c31c0db1388e9c23c4859e239824bdf29059c5a812c3ea501f3900000000:
      256'h4820a4a4c044b523a5c292556b0d89125df0a0a6da59a78b953571bf58d6d884;
        data[127] = 'd512 + 'hf89;
    end else begin
      compression = opcode_i[0] ?
      256'hb1d2c4905656d571f7ef0806f590be218c814f386ab117310a8d381800000000:
      256'h0637697e16c69aaf54c92a0a4338ba4318235f7ca65937afaf39e5387e06784b;
    end
  #1; endtask
  //09a09c09c989a09023b432e28000323f87c79a9008f0ff323225656e3326234fca889df080bc09a3bc54d2af4b23c26e32bb2af423e2a24c4f5233c599c7689e
  task automatic assigning_key();
    key[0:15] = { 32'h09a09c09, 32'hc989a090,
                  32'h23b432e2, 32'h8000323f,
                  32'h87c79a90, 32'h08f0ff32,
                  32'h3225656e, 32'h3326234f,
                  32'hca889df0, 32'h80bc09a3,
                  32'hbc54d2af, 32'h4b23c26e,
                  32'h32bb2af4, 32'h23e2a24c,
                  32'h4f5233c5, 32'h99c7689e };
  #1; endtask
  
  task automatic assigning_simple_key();
    key[0:15] = { 32'h0000000c, 32'h0000000d,
                  32'h0000000a, 32'h0000000b,
                  32'h00000008, 32'h00000009,
                  32'h00000090, 32'h00000080,
                  32'h000000f0, 32'h000000e0,
                  32'h000000d0, 32'h000000c0,
                  32'h00000c00, 32'h00000d00,
                  32'h00000a00, 32'h00000b0f };
  #1; endtask
  
  task automatic assigning_title(); #1
    case (opcode_i)
      0: begin mode = "sha 256: "; m = sha_256; end
      1: begin mode = "sha 244: "; m = sha_224; end
      2: begin mode = "HMAC 256: "; m = HMAC_256; end
      3: begin mode = "HMAC 224: "; m = HMAC_224; end
    endcase
  endtask
  
  task automatic running_tests(input [1:0] opcode);
    #1 opcode_i = opcode;assigning_title(); test_vec_1(); SendBlockData(1); 
    #1 opcode_i = opcode;assigning_title(); test_vec_2(); SendBlockData(1); 
    #1 opcode_i = opcode;assigning_title(); test_vec_3(); SendBlockData(2);
    #1 opcode_i = opcode;assigning_title(); test_vec_4(); SendBlockData(3);
    #1 opcode_i = opcode;assigning_title(); test_vec_5(); SendBlockData(6);
    #1 opcode_i = opcode;assigning_title(); test_vec_6(); SendBlockData(6);
    #1 opcode_i = opcode;assigning_title(); test_vec_7(); SendBlockData(8);
  endtask
  //////////////////////////////////////////////////////
  initial begin
    aresetn_i <= 0; #20
    aresetn_i <= 1;
    //////////////////////////////////////////////////////
//    assigning_simple_key();
    assigning_key();
    running_tests(0);
    running_tests(1);
    running_tests(2);
    running_tests(3);
  end
`endif `endif
endmodule
