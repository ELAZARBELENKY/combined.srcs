`timescale 1ns / 1ps
  //Address map
  localparam ID_ADDR   = 12'h000;
  localparam CFG_ADDR  = 12'h010;
  localparam CTL_ADDR  = 12'h020;
  localparam STS_ADDR  = 12'h030;
  localparam IE_ADDR   = 12'h040;
  localparam HASH_ADDR = 12'h100;
  localparam DIN_ADDR  = 12'h140;
  localparam KEY_ADDR  = 12'h150;
//  localparam SEED_ADDR = 12'h300;

module lw_sha_interface_control_logic #(
   parameter int FIQSHA_BUS_DATA_WIDTH = `FIQSHA_BUS,
   parameter int ARCH_SZ = `WORD_SIZE,
   parameter logic [31:0] ID_VAL = 32'h0)
   (
   input clk_i,
   input resetn_i,
   input wr_i,                                        // write from bus interface adapter
   output reg wr_ack_o,                               // write ackowledge to bus interface adapter
   input rd_i,                                        // read request from bus interface adapter
   input rd_ack_i,                                    // read ack from bus interface adapter
   input [11:0] waddr_i,                              // write address
   input [11:0] raddr_i,                              // read adress
   input [FIQSHA_BUS_DATA_WIDTH-1:0] wdata_i,         // write data
   output reg [FIQSHA_BUS_DATA_WIDTH-1:0] rdata_o,    // read data
   output reg read_valid_o,                           // read data validation strob
`ifdef HMACAUXKEY
   input [`KEY_SIZE-1:0] aux_key_i, // dedicated key port to protected secret input instead bus transaction.
`endif

   input [1:0] burst_type_i,
   output irq_o,
   input overflow,
  // native interface
   input [`WORD_SIZE-1:0] hash_i[7:0],
   input ready_i,
   output new_key_o,
   input core_ready_i,
   input done_i,
   input fault_inj_det_i,
   input key_ready_i,
   output logic key_valid_o,
   output logic [`WORD_SIZE-1:0] key_o,
   output [`WORD_SIZE-1:0] data_o,
   output start_o,
   output abort_o,
   output last_o,
   output [3:0] opcode_o,
   output logic valid_o,
   
   output dma_wr_req_o,
   output dma_rd_req_o,
   output reg slv_error_o,
   output core_reset_o
   );
  
  localparam byte BUS_DATA_IN_ARCH_SZ = (ARCH_SZ + FIQSHA_BUS_DATA_WIDTH - 1)/FIQSHA_BUS_DATA_WIDTH;
  logic first_word = 1;
  logic s64;
  logic hash_avliable = 1'b0;
  logic [31:0] id_reg = ID_VAL;
  logic [31:0] cfg_reg, ctl_reg, sts_reg, ie_reg, seed_reg;
  logic [`WORD_SIZE-1:0] din_reg;
  logic [8*`WORD_SIZE-1:0] hash_reg;
  assign slv_error_o = wr_i && (waddr_i == DIN_ADDR && !ready_i ||
                                waddr_i == KEY_ADDR && !key_ready_i);
  localparam HASH_SIZE = `WORD_SIZE*8;
  assign wr_ack_o = wr_i;
  always_ff @(posedge clk_i or negedge resetn_i) begin
    if (~resetn_i) begin
      cfg_reg <= '0;
      ctl_reg <= '0;
      sts_reg[3] <= 1'b0;
      ie_reg <= 32'h2;
      seed_reg <= '0;
    end else begin
      if (overflow) sts_reg[6] <= 1'b1;
      if (wr_i) begin
//        wr_ack_o = 1'b1;
        case (waddr_i)
          CFG_ADDR: begin
            cfg_reg[7:0] <= wdata_i[7:0];
            cfg_reg[31] <= wdata_i[31];
          end
          CTL_ADDR: begin
            ctl_reg[31:0] <= {29'h0, wdata_i[2:0]};
            valid_o <= wdata_i[0] && (core_ready_i);
          end
          STS_ADDR: begin
            if (wdata_i[6]) sts_reg[6] <= 1'b0;
            if (wdata_i[3]) sts_reg[3] <= 1'b0;
            if (wdata_i[0]) sts_reg[0] <= 1'b0;
//            if (wdata_i & 4'b0110 != '0) slv_error_o <= 1'b1; 
          end
          IE_ADDR: begin
            ie_reg <= {27'h0, wdata_i[6:0]};
          end
          DIN_ADDR: begin
            if (ready_i) begin
`ifdef CORE_ARCH_S64
              if (`FIQSHA_BUS == 32 && s64) begin
                if (first_word) begin
                  din_reg[`WORD_SIZE-1-:`WORD_SIZE] <= wdata_i << 32;
                end else begin
                  din_reg[`WORD_SIZE/2-1:0] <= wdata_i;
                end
                valid_o <= !first_word;
                first_word <= !first_word;
              end else begin
                din_reg <= wdata_i;
                valid_o <= 1'b1;
              end
`else `ifdef CORE_ARCH_S32
              din_reg <= wdata_i;
              valid_o <= 1'b1;
`endif `endif
            end else begin
              sts_reg[3] <= 1'b1;
//              slv_error_o <= 1'b1;
            end
          end
`ifndef HMACAUXKEY
          KEY_ADDR: begin
            if (key_ready_i) begin
`ifdef CORE_ARCH_S64
              if (`FIQSHA_BUS == 32 && s64) begin
                if (first_word) begin
                  key_o[`WORD_SIZE-1-:`WORD_SIZE] <= wdata_i << 32;
                end else begin
                  key_o[`WORD_SIZE/2-1:0] <= wdata_i;
                end
                key_valid_o <= !first_word;
                first_word <= !first_word;
              end else begin
                key_o <= wdata_i;
                key_valid_o <= 1'b1;
              end
`else `ifdef CORE_ARCH_S32
              key_o <= wdata_i;
              key_valid_o <= 1'b1;
`endif `endif
            end else begin
              sts_reg[3] <= 1'b1;
//              slv_error_o <= 1'b1;
            end
          end
`endif
          default:;
        endcase
        if (cfg_reg[31]) begin
          cfg_reg <= '0;
          ctl_reg <= '0;
          sts_reg[6] <= '0;
          sts_reg[3] <= '1;
          ie_reg <= 32'h2;
        end
      end else begin
//        slv_error_o <= 1'b0;
//        wr_ack_o = 1'b0;
        if (start_o) ctl_reg[0] <= 1'b0;
        if (done_i) ctl_reg[1] <= 1'b0;
        if (abort_o) ctl_reg[2] <= 1'b0;
        valid_o <= 0;
`ifndef HMACAUXKEY
        key_valid_o <= 0;
`endif
      end
    end
  end
  
  wire [$clog2(HASH_SIZE/8)-$clog2(FIQSHA_BUS_DATA_WIDTH/8)-1:0] hash_reg_word_rptr = 
    raddr_i[$clog2(HASH_SIZE/8)-1:$clog2(FIQSHA_BUS_DATA_WIDTH/8)];
  
  always_ff @(posedge clk_i or negedge resetn_i) begin
    if (!resetn_i || start_o) hash_avliable <= 1'b0;
    else if (done_i) hash_avliable <= 1'b1;
  end

  always_comb begin
    rdata_o = '0;
    read_valid_o = 1'b0;
    if (!resetn_i) begin
      rdata_o = 32'h0;
      read_valid_o = 1'b1;
    end else if (rd_i) begin
      case (raddr_i)
        CFG_ADDR: begin
          rdata_o = {1'b0, cfg_reg[30:0]};
          read_valid_o = 1'b1;
        end
        CTL_ADDR: begin
          rdata_o = {ctl_reg[31:3], 3'b0};
          read_valid_o = 1'b1;
        end
        STS_ADDR: begin
          rdata_o = sts_reg;
          read_valid_o = 1'b1;
        end
        IE_ADDR: begin
          rdata_o = ie_reg;
          read_valid_o = 1'b1;
        end
        default: begin
          if (raddr_i[11:$clog2(`WORD_SIZE)] === HASH_ADDR[11:$clog2(`WORD_SIZE)]) begin
            for (int i = 0; i < HASH_SIZE/FIQSHA_BUS_DATA_WIDTH; i++) begin
              if (i === hash_reg_word_rptr)
                rdata_o = hash_reg[i*FIQSHA_BUS_DATA_WIDTH +: FIQSHA_BUS_DATA_WIDTH];
            end
            read_valid_o = 1'b1;
          end
        end
      endcase
    end
  end

  typedef struct {
    logic [15:0] majorid;
    logic [15:0] minorid;
  } id_t;

  typedef struct {
    logic srst;
    logic hmacnewkey;
    logic [3:0] opcode;
  } cfg_t;

  typedef struct {
    logic abort;
    logic last;
    logic init;
  } ctl_t;

  typedef struct {
    logic overflow;
    logic faultinjdet;
    logic busy;
    logic derr;
`ifndef HMACAUXKEY
    logic rdyk;
`endif
    logic rdyd;
    logic avl;
  } sts_t;

  typedef struct {
    logic overflow;
    logic faultinjdetie;
    logic busyie;
    logic derrie;
`ifndef HMACAUXKEY
    logic rdykie;
`endif
    logic rdydie;
    logic avlie;
  } ie_t;
  
  id_t id;
  cfg_t cfg;
  ctl_t ctl;
  sts_t sts;
  ie_t ie;

//  always_comb begin
   assign id = '{majorid: id_reg[31:16],
                 minorid: id_reg[15:0]};

   assign cfg = '{srst: cfg_reg[31],
                  hmacnewkey: cfg_reg[4],
                  opcode: cfg_reg[3:0]};

   assign ctl = '{abort: ctl_reg[2],
                  last: ctl_reg[1],
                  init: ctl_reg[0]};

   assign sts = '{overflow: sts_reg[6],
                  faultinjdet: sts_reg[5],
                  busy: sts_reg[4],
                  derr: sts_reg[3],
`ifndef HMACAUXKEY
                  rdyk: sts_reg[2],
`endif
                  rdyd: sts_reg[1],
                  avl: sts_reg[0]};

    assign ie = '{overflow: ie_reg[6],
                  faultinjdetie: ie_reg[5],
                  busyie: ie_reg[4],
                  derrie: ie_reg[3],
`ifndef HMACAUXKEY
                  rdykie: ie_reg[2],
`endif
                  rdydie: ie_reg[1],
                  avlie: ie_reg[0]};
//  end

  assign hash_reg = {hash_i[7],hash_i[6],hash_i[5],hash_i[4],
                     hash_i[3],hash_i[2],hash_i[1],hash_i[0]};
  assign sts_reg[5:4] = {fault_inj_det_i, !core_ready_i};
  assign sts_reg[1:0] = {ready_i, done_i || hash_avliable};
  assign sts_reg[31:5] = '0;
  assign start_o = ctl.init;
  assign last_o = ctl.last;
  assign abort_o = ctl.abort;
  assign opcode_o = cfg.opcode;
  assign new_key_o = cfg.hmacnewkey;
  assign core_reset_o = !cfg.srst;
  assign data_o = din_reg;
  assign dma_wr_req_o = sts.rdyd;
  assign dma_rd_req_o = sts.avl;
`ifndef HMACAUXKEY
  assign sts_reg[2] = key_ready_i;
`else
  assign sts_reg[2] = 1'b0;
`endif

`ifdef CORE_ARCH_S64
  assign s64 = cfg.opcode[3]||cfg.opcode[2];
`else `ifdef CORE_ARCH_S32
  assign s64 = 1'b1;
`endif `endif
  assign irq_o =
     (sts.overflow & ie.overflow) |
     (sts.faultinjdet & ie.faultinjdetie) |
     (sts.busy & ie.busyie) |
     (sts.derr & ie.derrie) |
`ifndef HMACAUXKEY
     (sts.rdyk & ie.rdykie) |
`endif
     (sts.rdyd & ie.rdydie) |
     (sts.avl & ie.avlie);

`ifdef HMACAUXKEY
  
  localparam int max_ctr = `KEY_SIZE/`WORD_SIZE;
  localparam longint mask = {`KEY_SIZE%`WORD_SIZE{1'b1}}<<`WORD_SIZE-`KEY_SIZE%`WORD_SIZE;
`ifdef CORE_ARCH_S64
  localparam logic div_mask = `KEY_SIZE%`WORD_SIZE < `WORD_SIZE/2;
  localparam logic good_key = `KEY_SIZE <= 512;
  logic [`SAFE_CLOG2(`KEY_SIZE/`WORD_SIZE):0] ctr = 0;
`else `ifdef CORE_ARCH_S32
  logic [`SAFE_CLOG2(`KEY_SIZE/`WORD_SIZE)-1:0] ctr = 0;
`endif `endif
  logic [`SAFE_CLOG2(`KEY_SIZE)-1:0] ptr;
  logic key_zero;
  
`ifdef CORE_ARCH_S64
  assign ptr = `KEY_SIZE-(s64||good_key?0:`KEY_SIZE-512)-ctr*`WORD_SIZE/(s64?1:2)-1;
`else `ifdef CORE_ARCH_S32
  assign ptr = `KEY_SIZE-ctr*`WORD_SIZE-1;
`endif `endif

  always_ff @(posedge clk_i) begin
    key_valid_o <= key_ready_i;
    if (key_ready_i) begin
      if (key_zero) key_o <= '0;
`ifdef CORE_ARCH_S64
      else if (ctr == max_ctr*(s64?1:2)+(!s64&&!div_mask)) begin
        key_o <= (s64 ? aux_key_i[ptr-:`WORD_SIZE]:
        aux_key_i[ptr-:`WORD_SIZE/2]) & (mask >> (!s64&&div_mask?32:0));
`else `ifdef CORE_ARCH_S32
      else if (ctr == max_ctr) begin
        key_o <= aux_key_i[ptr-:`WORD_SIZE] & mask;
`endif `endif
        key_zero <= 1'b1;
      end else begin
        key_o <= (s64 ? aux_key_i[ptr-:`WORD_SIZE]:
                        aux_key_i[ptr-:`WORD_SIZE/2]);
        ctr <= ctr + 1;
      end
    end else if (start_o) begin
      key_zero <= 1'b0;
      ctr <= 0;
    end
  end
`endif
endmodule
